module wave_table_test(
					  input logic [12:0] ADDR,
					  output logic [15:0] SAMPLE
					  );
					  
always_comb begin

	case(ADDR)
		0: SAMPLE = 16'h0;
		1: SAMPLE = 16'h32;
		2: SAMPLE = 16'h64;
		3: SAMPLE = 16'h96;
		4: SAMPLE = 16'hc9;
		5: SAMPLE = 16'hfb;
		6: SAMPLE = 16'h12d;
		7: SAMPLE = 16'h15f;
		8: SAMPLE = 16'h192;
		9: SAMPLE = 16'h1c4;
		10: SAMPLE = 16'h1f6;
		11: SAMPLE = 16'h228;
		12: SAMPLE = 16'h25b;
		13: SAMPLE = 16'h28d;
		14: SAMPLE = 16'h2bf;
		15: SAMPLE = 16'h2f1;
		16: SAMPLE = 16'h324;
		17: SAMPLE = 16'h356;
		18: SAMPLE = 16'h388;
		19: SAMPLE = 16'h3ba;
		20: SAMPLE = 16'h3ed;
		21: SAMPLE = 16'h41f;
		22: SAMPLE = 16'h451;
		23: SAMPLE = 16'h483;
		24: SAMPLE = 16'h4b6;
		25: SAMPLE = 16'h4e8;
		26: SAMPLE = 16'h51a;
		27: SAMPLE = 16'h54c;
		28: SAMPLE = 16'h57f;
		29: SAMPLE = 16'h5b1;
		30: SAMPLE = 16'h5e3;
		31: SAMPLE = 16'h615;
		32: SAMPLE = 16'h647;
		33: SAMPLE = 16'h67a;
		34: SAMPLE = 16'h6ac;
		35: SAMPLE = 16'h6de;
		36: SAMPLE = 16'h710;
		37: SAMPLE = 16'h742;
		38: SAMPLE = 16'h775;
		39: SAMPLE = 16'h7a7;
		40: SAMPLE = 16'h7d9;
		41: SAMPLE = 16'h80b;
		42: SAMPLE = 16'h83d;
		43: SAMPLE = 16'h86f;
		44: SAMPLE = 16'h8a2;
		45: SAMPLE = 16'h8d4;
		46: SAMPLE = 16'h906;
		47: SAMPLE = 16'h938;
		48: SAMPLE = 16'h96a;
		49: SAMPLE = 16'h99c;
		50: SAMPLE = 16'h9ce;
		51: SAMPLE = 16'ha00;
		52: SAMPLE = 16'ha33;
		53: SAMPLE = 16'ha65;
		54: SAMPLE = 16'ha97;
		55: SAMPLE = 16'hac9;
		56: SAMPLE = 16'hafb;
		57: SAMPLE = 16'hb2d;
		58: SAMPLE = 16'hb5f;
		59: SAMPLE = 16'hb91;
		60: SAMPLE = 16'hbc3;
		61: SAMPLE = 16'hbf5;
		62: SAMPLE = 16'hc27;
		63: SAMPLE = 16'hc59;
		64: SAMPLE = 16'hc8b;
		65: SAMPLE = 16'hcbd;
		66: SAMPLE = 16'hcef;
		67: SAMPLE = 16'hd21;
		68: SAMPLE = 16'hd53;
		69: SAMPLE = 16'hd85;
		70: SAMPLE = 16'hdb7;
		71: SAMPLE = 16'hde9;
		72: SAMPLE = 16'he1b;
		73: SAMPLE = 16'he4d;
		74: SAMPLE = 16'he7f;
		75: SAMPLE = 16'heb1;
		76: SAMPLE = 16'hee3;
		77: SAMPLE = 16'hf15;
		78: SAMPLE = 16'hf47;
		79: SAMPLE = 16'hf79;
		80: SAMPLE = 16'hfab;
		81: SAMPLE = 16'hfdd;
		82: SAMPLE = 16'h100e;
		83: SAMPLE = 16'h1040;
		84: SAMPLE = 16'h1072;
		85: SAMPLE = 16'h10a4;
		86: SAMPLE = 16'h10d6;
		87: SAMPLE = 16'h1108;
		88: SAMPLE = 16'h1139;
		89: SAMPLE = 16'h116b;
		90: SAMPLE = 16'h119d;
		91: SAMPLE = 16'h11cf;
		92: SAMPLE = 16'h1201;
		93: SAMPLE = 16'h1232;
		94: SAMPLE = 16'h1264;
		95: SAMPLE = 16'h1296;
		96: SAMPLE = 16'h12c8;
		97: SAMPLE = 16'h12f9;
		98: SAMPLE = 16'h132b;
		99: SAMPLE = 16'h135d;
		100: SAMPLE = 16'h138e;
		101: SAMPLE = 16'h13c0;
		102: SAMPLE = 16'h13f2;
		103: SAMPLE = 16'h1423;
		104: SAMPLE = 16'h1455;
		105: SAMPLE = 16'h1487;
		106: SAMPLE = 16'h14b8;
		107: SAMPLE = 16'h14ea;
		108: SAMPLE = 16'h151b;
		109: SAMPLE = 16'h154d;
		110: SAMPLE = 16'h157f;
		111: SAMPLE = 16'h15b0;
		112: SAMPLE = 16'h15e2;
		113: SAMPLE = 16'h1613;
		114: SAMPLE = 16'h1645;
		115: SAMPLE = 16'h1676;
		116: SAMPLE = 16'h16a8;
		117: SAMPLE = 16'h16d9;
		118: SAMPLE = 16'h170a;
		119: SAMPLE = 16'h173c;
		120: SAMPLE = 16'h176d;
		121: SAMPLE = 16'h179f;
		122: SAMPLE = 16'h17d0;
		123: SAMPLE = 16'h1802;
		124: SAMPLE = 16'h1833;
		125: SAMPLE = 16'h1864;
		126: SAMPLE = 16'h1896;
		127: SAMPLE = 16'h18c7;
		128: SAMPLE = 16'h18f8;
		129: SAMPLE = 16'h192a;
		130: SAMPLE = 16'h195b;
		131: SAMPLE = 16'h198c;
		132: SAMPLE = 16'h19bd;
		133: SAMPLE = 16'h19ef;
		134: SAMPLE = 16'h1a20;
		135: SAMPLE = 16'h1a51;
		136: SAMPLE = 16'h1a82;
		137: SAMPLE = 16'h1ab3;
		138: SAMPLE = 16'h1ae4;
		139: SAMPLE = 16'h1b16;
		140: SAMPLE = 16'h1b47;
		141: SAMPLE = 16'h1b78;
		142: SAMPLE = 16'h1ba9;
		143: SAMPLE = 16'h1bda;
		144: SAMPLE = 16'h1c0b;
		145: SAMPLE = 16'h1c3c;
		146: SAMPLE = 16'h1c6d;
		147: SAMPLE = 16'h1c9e;
		148: SAMPLE = 16'h1ccf;
		149: SAMPLE = 16'h1d00;
		150: SAMPLE = 16'h1d31;
		151: SAMPLE = 16'h1d62;
		152: SAMPLE = 16'h1d93;
		153: SAMPLE = 16'h1dc4;
		154: SAMPLE = 16'h1df5;
		155: SAMPLE = 16'h1e25;
		156: SAMPLE = 16'h1e56;
		157: SAMPLE = 16'h1e87;
		158: SAMPLE = 16'h1eb8;
		159: SAMPLE = 16'h1ee9;
		160: SAMPLE = 16'h1f19;
		161: SAMPLE = 16'h1f4a;
		162: SAMPLE = 16'h1f7b;
		163: SAMPLE = 16'h1fac;
		164: SAMPLE = 16'h1fdc;
		165: SAMPLE = 16'h200d;
		166: SAMPLE = 16'h203e;
		167: SAMPLE = 16'h206e;
		168: SAMPLE = 16'h209f;
		169: SAMPLE = 16'h20d0;
		170: SAMPLE = 16'h2100;
		171: SAMPLE = 16'h2131;
		172: SAMPLE = 16'h2161;
		173: SAMPLE = 16'h2192;
		174: SAMPLE = 16'h21c2;
		175: SAMPLE = 16'h21f3;
		176: SAMPLE = 16'h2223;
		177: SAMPLE = 16'h2254;
		178: SAMPLE = 16'h2284;
		179: SAMPLE = 16'h22b4;
		180: SAMPLE = 16'h22e5;
		181: SAMPLE = 16'h2315;
		182: SAMPLE = 16'h2345;
		183: SAMPLE = 16'h2376;
		184: SAMPLE = 16'h23a6;
		185: SAMPLE = 16'h23d6;
		186: SAMPLE = 16'h2407;
		187: SAMPLE = 16'h2437;
		188: SAMPLE = 16'h2467;
		189: SAMPLE = 16'h2497;
		190: SAMPLE = 16'h24c7;
		191: SAMPLE = 16'h24f7;
		192: SAMPLE = 16'h2528;
		193: SAMPLE = 16'h2558;
		194: SAMPLE = 16'h2588;
		195: SAMPLE = 16'h25b8;
		196: SAMPLE = 16'h25e8;
		197: SAMPLE = 16'h2618;
		198: SAMPLE = 16'h2648;
		199: SAMPLE = 16'h2678;
		200: SAMPLE = 16'h26a8;
		201: SAMPLE = 16'h26d8;
		202: SAMPLE = 16'h2707;
		203: SAMPLE = 16'h2737;
		204: SAMPLE = 16'h2767;
		205: SAMPLE = 16'h2797;
		206: SAMPLE = 16'h27c7;
		207: SAMPLE = 16'h27f6;
		208: SAMPLE = 16'h2826;
		209: SAMPLE = 16'h2856;
		210: SAMPLE = 16'h2886;
		211: SAMPLE = 16'h28b5;
		212: SAMPLE = 16'h28e5;
		213: SAMPLE = 16'h2915;
		214: SAMPLE = 16'h2944;
		215: SAMPLE = 16'h2974;
		216: SAMPLE = 16'h29a3;
		217: SAMPLE = 16'h29d3;
		218: SAMPLE = 16'h2a02;
		219: SAMPLE = 16'h2a32;
		220: SAMPLE = 16'h2a61;
		221: SAMPLE = 16'h2a91;
		222: SAMPLE = 16'h2ac0;
		223: SAMPLE = 16'h2aef;
		224: SAMPLE = 16'h2b1f;
		225: SAMPLE = 16'h2b4e;
		226: SAMPLE = 16'h2b7d;
		227: SAMPLE = 16'h2bad;
		228: SAMPLE = 16'h2bdc;
		229: SAMPLE = 16'h2c0b;
		230: SAMPLE = 16'h2c3a;
		231: SAMPLE = 16'h2c69;
		232: SAMPLE = 16'h2c98;
		233: SAMPLE = 16'h2cc8;
		234: SAMPLE = 16'h2cf7;
		235: SAMPLE = 16'h2d26;
		236: SAMPLE = 16'h2d55;
		237: SAMPLE = 16'h2d84;
		238: SAMPLE = 16'h2db3;
		239: SAMPLE = 16'h2de2;
		240: SAMPLE = 16'h2e11;
		241: SAMPLE = 16'h2e3f;
		242: SAMPLE = 16'h2e6e;
		243: SAMPLE = 16'h2e9d;
		244: SAMPLE = 16'h2ecc;
		245: SAMPLE = 16'h2efb;
		246: SAMPLE = 16'h2f29;
		247: SAMPLE = 16'h2f58;
		248: SAMPLE = 16'h2f87;
		249: SAMPLE = 16'h2fb5;
		250: SAMPLE = 16'h2fe4;
		251: SAMPLE = 16'h3013;
		252: SAMPLE = 16'h3041;
		253: SAMPLE = 16'h3070;
		254: SAMPLE = 16'h309e;
		255: SAMPLE = 16'h30cd;
		256: SAMPLE = 16'h30fb;
		257: SAMPLE = 16'h312a;
		258: SAMPLE = 16'h3158;
		259: SAMPLE = 16'h3186;
		260: SAMPLE = 16'h31b5;
		261: SAMPLE = 16'h31e3;
		262: SAMPLE = 16'h3211;
		263: SAMPLE = 16'h3240;
		264: SAMPLE = 16'h326e;
		265: SAMPLE = 16'h329c;
		266: SAMPLE = 16'h32ca;
		267: SAMPLE = 16'h32f8;
		268: SAMPLE = 16'h3326;
		269: SAMPLE = 16'h3354;
		270: SAMPLE = 16'h3382;
		271: SAMPLE = 16'h33b0;
		272: SAMPLE = 16'h33de;
		273: SAMPLE = 16'h340c;
		274: SAMPLE = 16'h343a;
		275: SAMPLE = 16'h3468;
		276: SAMPLE = 16'h3496;
		277: SAMPLE = 16'h34c4;
		278: SAMPLE = 16'h34f2;
		279: SAMPLE = 16'h351f;
		280: SAMPLE = 16'h354d;
		281: SAMPLE = 16'h357b;
		282: SAMPLE = 16'h35a8;
		283: SAMPLE = 16'h35d6;
		284: SAMPLE = 16'h3604;
		285: SAMPLE = 16'h3631;
		286: SAMPLE = 16'h365f;
		287: SAMPLE = 16'h368c;
		288: SAMPLE = 16'h36ba;
		289: SAMPLE = 16'h36e7;
		290: SAMPLE = 16'h3714;
		291: SAMPLE = 16'h3742;
		292: SAMPLE = 16'h376f;
		293: SAMPLE = 16'h379c;
		294: SAMPLE = 16'h37ca;
		295: SAMPLE = 16'h37f7;
		296: SAMPLE = 16'h3824;
		297: SAMPLE = 16'h3851;
		298: SAMPLE = 16'h387e;
		299: SAMPLE = 16'h38ab;
		300: SAMPLE = 16'h38d8;
		301: SAMPLE = 16'h3906;
		302: SAMPLE = 16'h3932;
		303: SAMPLE = 16'h395f;
		304: SAMPLE = 16'h398c;
		305: SAMPLE = 16'h39b9;
		306: SAMPLE = 16'h39e6;
		307: SAMPLE = 16'h3a13;
		308: SAMPLE = 16'h3a40;
		309: SAMPLE = 16'h3a6c;
		310: SAMPLE = 16'h3a99;
		311: SAMPLE = 16'h3ac6;
		312: SAMPLE = 16'h3af2;
		313: SAMPLE = 16'h3b1f;
		314: SAMPLE = 16'h3b4c;
		315: SAMPLE = 16'h3b78;
		316: SAMPLE = 16'h3ba5;
		317: SAMPLE = 16'h3bd1;
		318: SAMPLE = 16'h3bfd;
		319: SAMPLE = 16'h3c2a;
		320: SAMPLE = 16'h3c56;
		321: SAMPLE = 16'h3c83;
		322: SAMPLE = 16'h3caf;
		323: SAMPLE = 16'h3cdb;
		324: SAMPLE = 16'h3d07;
		325: SAMPLE = 16'h3d33;
		326: SAMPLE = 16'h3d60;
		327: SAMPLE = 16'h3d8c;
		328: SAMPLE = 16'h3db8;
		329: SAMPLE = 16'h3de4;
		330: SAMPLE = 16'h3e10;
		331: SAMPLE = 16'h3e3c;
		332: SAMPLE = 16'h3e68;
		333: SAMPLE = 16'h3e93;
		334: SAMPLE = 16'h3ebf;
		335: SAMPLE = 16'h3eeb;
		336: SAMPLE = 16'h3f17;
		337: SAMPLE = 16'h3f43;
		338: SAMPLE = 16'h3f6e;
		339: SAMPLE = 16'h3f9a;
		340: SAMPLE = 16'h3fc5;
		341: SAMPLE = 16'h3ff1;
		342: SAMPLE = 16'h401d;
		343: SAMPLE = 16'h4048;
		344: SAMPLE = 16'h4073;
		345: SAMPLE = 16'h409f;
		346: SAMPLE = 16'h40ca;
		347: SAMPLE = 16'h40f6;
		348: SAMPLE = 16'h4121;
		349: SAMPLE = 16'h414c;
		350: SAMPLE = 16'h4177;
		351: SAMPLE = 16'h41a2;
		352: SAMPLE = 16'h41ce;
		353: SAMPLE = 16'h41f9;
		354: SAMPLE = 16'h4224;
		355: SAMPLE = 16'h424f;
		356: SAMPLE = 16'h427a;
		357: SAMPLE = 16'h42a5;
		358: SAMPLE = 16'h42d0;
		359: SAMPLE = 16'h42fa;
		360: SAMPLE = 16'h4325;
		361: SAMPLE = 16'h4350;
		362: SAMPLE = 16'h437b;
		363: SAMPLE = 16'h43a5;
		364: SAMPLE = 16'h43d0;
		365: SAMPLE = 16'h43fb;
		366: SAMPLE = 16'h4425;
		367: SAMPLE = 16'h4450;
		368: SAMPLE = 16'h447a;
		369: SAMPLE = 16'h44a5;
		370: SAMPLE = 16'h44cf;
		371: SAMPLE = 16'h44fa;
		372: SAMPLE = 16'h4524;
		373: SAMPLE = 16'h454e;
		374: SAMPLE = 16'h4578;
		375: SAMPLE = 16'h45a3;
		376: SAMPLE = 16'h45cd;
		377: SAMPLE = 16'h45f7;
		378: SAMPLE = 16'h4621;
		379: SAMPLE = 16'h464b;
		380: SAMPLE = 16'h4675;
		381: SAMPLE = 16'h469f;
		382: SAMPLE = 16'h46c9;
		383: SAMPLE = 16'h46f3;
		384: SAMPLE = 16'h471c;
		385: SAMPLE = 16'h4746;
		386: SAMPLE = 16'h4770;
		387: SAMPLE = 16'h479a;
		388: SAMPLE = 16'h47c3;
		389: SAMPLE = 16'h47ed;
		390: SAMPLE = 16'h4816;
		391: SAMPLE = 16'h4840;
		392: SAMPLE = 16'h4869;
		393: SAMPLE = 16'h4893;
		394: SAMPLE = 16'h48bc;
		395: SAMPLE = 16'h48e6;
		396: SAMPLE = 16'h490f;
		397: SAMPLE = 16'h4938;
		398: SAMPLE = 16'h4961;
		399: SAMPLE = 16'h498a;
		400: SAMPLE = 16'h49b4;
		401: SAMPLE = 16'h49dd;
		402: SAMPLE = 16'h4a06;
		403: SAMPLE = 16'h4a2f;
		404: SAMPLE = 16'h4a58;
		405: SAMPLE = 16'h4a81;
		406: SAMPLE = 16'h4aa9;
		407: SAMPLE = 16'h4ad2;
		408: SAMPLE = 16'h4afb;
		409: SAMPLE = 16'h4b24;
		410: SAMPLE = 16'h4b4c;
		411: SAMPLE = 16'h4b75;
		412: SAMPLE = 16'h4b9e;
		413: SAMPLE = 16'h4bc6;
		414: SAMPLE = 16'h4bef;
		415: SAMPLE = 16'h4c17;
		416: SAMPLE = 16'h4c3f;
		417: SAMPLE = 16'h4c68;
		418: SAMPLE = 16'h4c90;
		419: SAMPLE = 16'h4cb8;
		420: SAMPLE = 16'h4ce1;
		421: SAMPLE = 16'h4d09;
		422: SAMPLE = 16'h4d31;
		423: SAMPLE = 16'h4d59;
		424: SAMPLE = 16'h4d81;
		425: SAMPLE = 16'h4da9;
		426: SAMPLE = 16'h4dd1;
		427: SAMPLE = 16'h4df9;
		428: SAMPLE = 16'h4e21;
		429: SAMPLE = 16'h4e48;
		430: SAMPLE = 16'h4e70;
		431: SAMPLE = 16'h4e98;
		432: SAMPLE = 16'h4ebf;
		433: SAMPLE = 16'h4ee7;
		434: SAMPLE = 16'h4f0f;
		435: SAMPLE = 16'h4f36;
		436: SAMPLE = 16'h4f5e;
		437: SAMPLE = 16'h4f85;
		438: SAMPLE = 16'h4fac;
		439: SAMPLE = 16'h4fd4;
		440: SAMPLE = 16'h4ffb;
		441: SAMPLE = 16'h5022;
		442: SAMPLE = 16'h5049;
		443: SAMPLE = 16'h5070;
		444: SAMPLE = 16'h5097;
		445: SAMPLE = 16'h50bf;
		446: SAMPLE = 16'h50e5;
		447: SAMPLE = 16'h510c;
		448: SAMPLE = 16'h5133;
		449: SAMPLE = 16'h515a;
		450: SAMPLE = 16'h5181;
		451: SAMPLE = 16'h51a8;
		452: SAMPLE = 16'h51ce;
		453: SAMPLE = 16'h51f5;
		454: SAMPLE = 16'h521c;
		455: SAMPLE = 16'h5242;
		456: SAMPLE = 16'h5269;
		457: SAMPLE = 16'h528f;
		458: SAMPLE = 16'h52b5;
		459: SAMPLE = 16'h52dc;
		460: SAMPLE = 16'h5302;
		461: SAMPLE = 16'h5328;
		462: SAMPLE = 16'h534e;
		463: SAMPLE = 16'h5375;
		464: SAMPLE = 16'h539b;
		465: SAMPLE = 16'h53c1;
		466: SAMPLE = 16'h53e7;
		467: SAMPLE = 16'h540d;
		468: SAMPLE = 16'h5433;
		469: SAMPLE = 16'h5458;
		470: SAMPLE = 16'h547e;
		471: SAMPLE = 16'h54a4;
		472: SAMPLE = 16'h54ca;
		473: SAMPLE = 16'h54ef;
		474: SAMPLE = 16'h5515;
		475: SAMPLE = 16'h553a;
		476: SAMPLE = 16'h5560;
		477: SAMPLE = 16'h5585;
		478: SAMPLE = 16'h55ab;
		479: SAMPLE = 16'h55d0;
		480: SAMPLE = 16'h55f5;
		481: SAMPLE = 16'h561a;
		482: SAMPLE = 16'h5640;
		483: SAMPLE = 16'h5665;
		484: SAMPLE = 16'h568a;
		485: SAMPLE = 16'h56af;
		486: SAMPLE = 16'h56d4;
		487: SAMPLE = 16'h56f9;
		488: SAMPLE = 16'h571d;
		489: SAMPLE = 16'h5742;
		490: SAMPLE = 16'h5767;
		491: SAMPLE = 16'h578c;
		492: SAMPLE = 16'h57b0;
		493: SAMPLE = 16'h57d5;
		494: SAMPLE = 16'h57f9;
		495: SAMPLE = 16'h581e;
		496: SAMPLE = 16'h5842;
		497: SAMPLE = 16'h5867;
		498: SAMPLE = 16'h588b;
		499: SAMPLE = 16'h58af;
		500: SAMPLE = 16'h58d4;
		501: SAMPLE = 16'h58f8;
		502: SAMPLE = 16'h591c;
		503: SAMPLE = 16'h5940;
		504: SAMPLE = 16'h5964;
		505: SAMPLE = 16'h5988;
		506: SAMPLE = 16'h59ac;
		507: SAMPLE = 16'h59d0;
		508: SAMPLE = 16'h59f3;
		509: SAMPLE = 16'h5a17;
		510: SAMPLE = 16'h5a3b;
		511: SAMPLE = 16'h5a5e;
		512: SAMPLE = 16'h5a82;
		513: SAMPLE = 16'h5aa5;
		514: SAMPLE = 16'h5ac9;
		515: SAMPLE = 16'h5aec;
		516: SAMPLE = 16'h5b10;
		517: SAMPLE = 16'h5b33;
		518: SAMPLE = 16'h5b56;
		519: SAMPLE = 16'h5b79;
		520: SAMPLE = 16'h5b9d;
		521: SAMPLE = 16'h5bc0;
		522: SAMPLE = 16'h5be3;
		523: SAMPLE = 16'h5c06;
		524: SAMPLE = 16'h5c29;
		525: SAMPLE = 16'h5c4b;
		526: SAMPLE = 16'h5c6e;
		527: SAMPLE = 16'h5c91;
		528: SAMPLE = 16'h5cb4;
		529: SAMPLE = 16'h5cd6;
		530: SAMPLE = 16'h5cf9;
		531: SAMPLE = 16'h5d1b;
		532: SAMPLE = 16'h5d3e;
		533: SAMPLE = 16'h5d60;
		534: SAMPLE = 16'h5d83;
		535: SAMPLE = 16'h5da5;
		536: SAMPLE = 16'h5dc7;
		537: SAMPLE = 16'h5de9;
		538: SAMPLE = 16'h5e0b;
		539: SAMPLE = 16'h5e2d;
		540: SAMPLE = 16'h5e50;
		541: SAMPLE = 16'h5e71;
		542: SAMPLE = 16'h5e93;
		543: SAMPLE = 16'h5eb5;
		544: SAMPLE = 16'h5ed7;
		545: SAMPLE = 16'h5ef9;
		546: SAMPLE = 16'h5f1a;
		547: SAMPLE = 16'h5f3c;
		548: SAMPLE = 16'h5f5e;
		549: SAMPLE = 16'h5f7f;
		550: SAMPLE = 16'h5fa0;
		551: SAMPLE = 16'h5fc2;
		552: SAMPLE = 16'h5fe3;
		553: SAMPLE = 16'h6004;
		554: SAMPLE = 16'h6026;
		555: SAMPLE = 16'h6047;
		556: SAMPLE = 16'h6068;
		557: SAMPLE = 16'h6089;
		558: SAMPLE = 16'h60aa;
		559: SAMPLE = 16'h60cb;
		560: SAMPLE = 16'h60ec;
		561: SAMPLE = 16'h610d;
		562: SAMPLE = 16'h612d;
		563: SAMPLE = 16'h614e;
		564: SAMPLE = 16'h616f;
		565: SAMPLE = 16'h618f;
		566: SAMPLE = 16'h61b0;
		567: SAMPLE = 16'h61d0;
		568: SAMPLE = 16'h61f1;
		569: SAMPLE = 16'h6211;
		570: SAMPLE = 16'h6231;
		571: SAMPLE = 16'h6251;
		572: SAMPLE = 16'h6271;
		573: SAMPLE = 16'h6292;
		574: SAMPLE = 16'h62b2;
		575: SAMPLE = 16'h62d2;
		576: SAMPLE = 16'h62f2;
		577: SAMPLE = 16'h6311;
		578: SAMPLE = 16'h6331;
		579: SAMPLE = 16'h6351;
		580: SAMPLE = 16'h6371;
		581: SAMPLE = 16'h6390;
		582: SAMPLE = 16'h63b0;
		583: SAMPLE = 16'h63cf;
		584: SAMPLE = 16'h63ef;
		585: SAMPLE = 16'h640e;
		586: SAMPLE = 16'h642d;
		587: SAMPLE = 16'h644d;
		588: SAMPLE = 16'h646c;
		589: SAMPLE = 16'h648b;
		590: SAMPLE = 16'h64aa;
		591: SAMPLE = 16'h64c9;
		592: SAMPLE = 16'h64e8;
		593: SAMPLE = 16'h6507;
		594: SAMPLE = 16'h6526;
		595: SAMPLE = 16'h6545;
		596: SAMPLE = 16'h6563;
		597: SAMPLE = 16'h6582;
		598: SAMPLE = 16'h65a0;
		599: SAMPLE = 16'h65bf;
		600: SAMPLE = 16'h65dd;
		601: SAMPLE = 16'h65fc;
		602: SAMPLE = 16'h661a;
		603: SAMPLE = 16'h6639;
		604: SAMPLE = 16'h6657;
		605: SAMPLE = 16'h6675;
		606: SAMPLE = 16'h6693;
		607: SAMPLE = 16'h66b1;
		608: SAMPLE = 16'h66cf;
		609: SAMPLE = 16'h66ed;
		610: SAMPLE = 16'h670b;
		611: SAMPLE = 16'h6729;
		612: SAMPLE = 16'h6746;
		613: SAMPLE = 16'h6764;
		614: SAMPLE = 16'h6782;
		615: SAMPLE = 16'h679f;
		616: SAMPLE = 16'h67bd;
		617: SAMPLE = 16'h67da;
		618: SAMPLE = 16'h67f7;
		619: SAMPLE = 16'h6815;
		620: SAMPLE = 16'h6832;
		621: SAMPLE = 16'h684f;
		622: SAMPLE = 16'h686c;
		623: SAMPLE = 16'h6889;
		624: SAMPLE = 16'h68a6;
		625: SAMPLE = 16'h68c3;
		626: SAMPLE = 16'h68e0;
		627: SAMPLE = 16'h68fd;
		628: SAMPLE = 16'h6919;
		629: SAMPLE = 16'h6936;
		630: SAMPLE = 16'h6953;
		631: SAMPLE = 16'h696f;
		632: SAMPLE = 16'h698c;
		633: SAMPLE = 16'h69a8;
		634: SAMPLE = 16'h69c4;
		635: SAMPLE = 16'h69e1;
		636: SAMPLE = 16'h69fd;
		637: SAMPLE = 16'h6a19;
		638: SAMPLE = 16'h6a35;
		639: SAMPLE = 16'h6a51;
		640: SAMPLE = 16'h6a6d;
		641: SAMPLE = 16'h6a89;
		642: SAMPLE = 16'h6aa5;
		643: SAMPLE = 16'h6ac1;
		644: SAMPLE = 16'h6adc;
		645: SAMPLE = 16'h6af8;
		646: SAMPLE = 16'h6b13;
		647: SAMPLE = 16'h6b2f;
		648: SAMPLE = 16'h6b4a;
		649: SAMPLE = 16'h6b66;
		650: SAMPLE = 16'h6b81;
		651: SAMPLE = 16'h6b9c;
		652: SAMPLE = 16'h6bb8;
		653: SAMPLE = 16'h6bd3;
		654: SAMPLE = 16'h6bee;
		655: SAMPLE = 16'h6c09;
		656: SAMPLE = 16'h6c24;
		657: SAMPLE = 16'h6c3f;
		658: SAMPLE = 16'h6c59;
		659: SAMPLE = 16'h6c74;
		660: SAMPLE = 16'h6c8f;
		661: SAMPLE = 16'h6ca9;
		662: SAMPLE = 16'h6cc4;
		663: SAMPLE = 16'h6cde;
		664: SAMPLE = 16'h6cf9;
		665: SAMPLE = 16'h6d13;
		666: SAMPLE = 16'h6d2d;
		667: SAMPLE = 16'h6d48;
		668: SAMPLE = 16'h6d62;
		669: SAMPLE = 16'h6d7c;
		670: SAMPLE = 16'h6d96;
		671: SAMPLE = 16'h6db0;
		672: SAMPLE = 16'h6dca;
		673: SAMPLE = 16'h6de3;
		674: SAMPLE = 16'h6dfd;
		675: SAMPLE = 16'h6e17;
		676: SAMPLE = 16'h6e30;
		677: SAMPLE = 16'h6e4a;
		678: SAMPLE = 16'h6e63;
		679: SAMPLE = 16'h6e7d;
		680: SAMPLE = 16'h6e96;
		681: SAMPLE = 16'h6eaf;
		682: SAMPLE = 16'h6ec9;
		683: SAMPLE = 16'h6ee2;
		684: SAMPLE = 16'h6efb;
		685: SAMPLE = 16'h6f14;
		686: SAMPLE = 16'h6f2d;
		687: SAMPLE = 16'h6f46;
		688: SAMPLE = 16'h6f5f;
		689: SAMPLE = 16'h6f77;
		690: SAMPLE = 16'h6f90;
		691: SAMPLE = 16'h6fa9;
		692: SAMPLE = 16'h6fc1;
		693: SAMPLE = 16'h6fda;
		694: SAMPLE = 16'h6ff2;
		695: SAMPLE = 16'h700a;
		696: SAMPLE = 16'h7023;
		697: SAMPLE = 16'h703b;
		698: SAMPLE = 16'h7053;
		699: SAMPLE = 16'h706b;
		700: SAMPLE = 16'h7083;
		701: SAMPLE = 16'h709b;
		702: SAMPLE = 16'h70b3;
		703: SAMPLE = 16'h70cb;
		704: SAMPLE = 16'h70e2;
		705: SAMPLE = 16'h70fa;
		706: SAMPLE = 16'h7112;
		707: SAMPLE = 16'h7129;
		708: SAMPLE = 16'h7141;
		709: SAMPLE = 16'h7158;
		710: SAMPLE = 16'h716f;
		711: SAMPLE = 16'h7186;
		712: SAMPLE = 16'h719e;
		713: SAMPLE = 16'h71b5;
		714: SAMPLE = 16'h71cc;
		715: SAMPLE = 16'h71e3;
		716: SAMPLE = 16'h71fa;
		717: SAMPLE = 16'h7211;
		718: SAMPLE = 16'h7227;
		719: SAMPLE = 16'h723e;
		720: SAMPLE = 16'h7255;
		721: SAMPLE = 16'h726b;
		722: SAMPLE = 16'h7282;
		723: SAMPLE = 16'h7298;
		724: SAMPLE = 16'h72af;
		725: SAMPLE = 16'h72c5;
		726: SAMPLE = 16'h72db;
		727: SAMPLE = 16'h72f1;
		728: SAMPLE = 16'h7307;
		729: SAMPLE = 16'h731d;
		730: SAMPLE = 16'h7333;
		731: SAMPLE = 16'h7349;
		732: SAMPLE = 16'h735f;
		733: SAMPLE = 16'h7375;
		734: SAMPLE = 16'h738a;
		735: SAMPLE = 16'h73a0;
		736: SAMPLE = 16'h73b5;
		737: SAMPLE = 16'h73cb;
		738: SAMPLE = 16'h73e0;
		739: SAMPLE = 16'h73f6;
		740: SAMPLE = 16'h740b;
		741: SAMPLE = 16'h7420;
		742: SAMPLE = 16'h7435;
		743: SAMPLE = 16'h744a;
		744: SAMPLE = 16'h745f;
		745: SAMPLE = 16'h7474;
		746: SAMPLE = 16'h7489;
		747: SAMPLE = 16'h749e;
		748: SAMPLE = 16'h74b2;
		749: SAMPLE = 16'h74c7;
		750: SAMPLE = 16'h74db;
		751: SAMPLE = 16'h74f0;
		752: SAMPLE = 16'h7504;
		753: SAMPLE = 16'h7519;
		754: SAMPLE = 16'h752d;
		755: SAMPLE = 16'h7541;
		756: SAMPLE = 16'h7555;
		757: SAMPLE = 16'h7569;
		758: SAMPLE = 16'h757d;
		759: SAMPLE = 16'h7591;
		760: SAMPLE = 16'h75a5;
		761: SAMPLE = 16'h75b9;
		762: SAMPLE = 16'h75cc;
		763: SAMPLE = 16'h75e0;
		764: SAMPLE = 16'h75f4;
		765: SAMPLE = 16'h7607;
		766: SAMPLE = 16'h761b;
		767: SAMPLE = 16'h762e;
		768: SAMPLE = 16'h7641;
		769: SAMPLE = 16'h7654;
		770: SAMPLE = 16'h7668;
		771: SAMPLE = 16'h767b;
		772: SAMPLE = 16'h768e;
		773: SAMPLE = 16'h76a0;
		774: SAMPLE = 16'h76b3;
		775: SAMPLE = 16'h76c6;
		776: SAMPLE = 16'h76d9;
		777: SAMPLE = 16'h76eb;
		778: SAMPLE = 16'h76fe;
		779: SAMPLE = 16'h7710;
		780: SAMPLE = 16'h7723;
		781: SAMPLE = 16'h7735;
		782: SAMPLE = 16'h7747;
		783: SAMPLE = 16'h775a;
		784: SAMPLE = 16'h776c;
		785: SAMPLE = 16'h777e;
		786: SAMPLE = 16'h7790;
		787: SAMPLE = 16'h77a2;
		788: SAMPLE = 16'h77b4;
		789: SAMPLE = 16'h77c5;
		790: SAMPLE = 16'h77d7;
		791: SAMPLE = 16'h77e9;
		792: SAMPLE = 16'h77fa;
		793: SAMPLE = 16'h780c;
		794: SAMPLE = 16'h781d;
		795: SAMPLE = 16'h782e;
		796: SAMPLE = 16'h7840;
		797: SAMPLE = 16'h7851;
		798: SAMPLE = 16'h7862;
		799: SAMPLE = 16'h7873;
		800: SAMPLE = 16'h7884;
		801: SAMPLE = 16'h7895;
		802: SAMPLE = 16'h78a6;
		803: SAMPLE = 16'h78b6;
		804: SAMPLE = 16'h78c7;
		805: SAMPLE = 16'h78d8;
		806: SAMPLE = 16'h78e8;
		807: SAMPLE = 16'h78f9;
		808: SAMPLE = 16'h7909;
		809: SAMPLE = 16'h7919;
		810: SAMPLE = 16'h792a;
		811: SAMPLE = 16'h793a;
		812: SAMPLE = 16'h794a;
		813: SAMPLE = 16'h795a;
		814: SAMPLE = 16'h796a;
		815: SAMPLE = 16'h797a;
		816: SAMPLE = 16'h798a;
		817: SAMPLE = 16'h7999;
		818: SAMPLE = 16'h79a9;
		819: SAMPLE = 16'h79b9;
		820: SAMPLE = 16'h79c8;
		821: SAMPLE = 16'h79d8;
		822: SAMPLE = 16'h79e7;
		823: SAMPLE = 16'h79f6;
		824: SAMPLE = 16'h7a05;
		825: SAMPLE = 16'h7a15;
		826: SAMPLE = 16'h7a24;
		827: SAMPLE = 16'h7a33;
		828: SAMPLE = 16'h7a42;
		829: SAMPLE = 16'h7a50;
		830: SAMPLE = 16'h7a5f;
		831: SAMPLE = 16'h7a6e;
		832: SAMPLE = 16'h7a7d;
		833: SAMPLE = 16'h7a8b;
		834: SAMPLE = 16'h7a9a;
		835: SAMPLE = 16'h7aa8;
		836: SAMPLE = 16'h7ab6;
		837: SAMPLE = 16'h7ac5;
		838: SAMPLE = 16'h7ad3;
		839: SAMPLE = 16'h7ae1;
		840: SAMPLE = 16'h7aef;
		841: SAMPLE = 16'h7afd;
		842: SAMPLE = 16'h7b0b;
		843: SAMPLE = 16'h7b19;
		844: SAMPLE = 16'h7b26;
		845: SAMPLE = 16'h7b34;
		846: SAMPLE = 16'h7b42;
		847: SAMPLE = 16'h7b4f;
		848: SAMPLE = 16'h7b5d;
		849: SAMPLE = 16'h7b6a;
		850: SAMPLE = 16'h7b77;
		851: SAMPLE = 16'h7b84;
		852: SAMPLE = 16'h7b92;
		853: SAMPLE = 16'h7b9f;
		854: SAMPLE = 16'h7bac;
		855: SAMPLE = 16'h7bb9;
		856: SAMPLE = 16'h7bc5;
		857: SAMPLE = 16'h7bd2;
		858: SAMPLE = 16'h7bdf;
		859: SAMPLE = 16'h7beb;
		860: SAMPLE = 16'h7bf8;
		861: SAMPLE = 16'h7c05;
		862: SAMPLE = 16'h7c11;
		863: SAMPLE = 16'h7c1d;
		864: SAMPLE = 16'h7c29;
		865: SAMPLE = 16'h7c36;
		866: SAMPLE = 16'h7c42;
		867: SAMPLE = 16'h7c4e;
		868: SAMPLE = 16'h7c5a;
		869: SAMPLE = 16'h7c66;
		870: SAMPLE = 16'h7c71;
		871: SAMPLE = 16'h7c7d;
		872: SAMPLE = 16'h7c89;
		873: SAMPLE = 16'h7c94;
		874: SAMPLE = 16'h7ca0;
		875: SAMPLE = 16'h7cab;
		876: SAMPLE = 16'h7cb7;
		877: SAMPLE = 16'h7cc2;
		878: SAMPLE = 16'h7ccd;
		879: SAMPLE = 16'h7cd8;
		880: SAMPLE = 16'h7ce3;
		881: SAMPLE = 16'h7cee;
		882: SAMPLE = 16'h7cf9;
		883: SAMPLE = 16'h7d04;
		884: SAMPLE = 16'h7d0f;
		885: SAMPLE = 16'h7d19;
		886: SAMPLE = 16'h7d24;
		887: SAMPLE = 16'h7d2f;
		888: SAMPLE = 16'h7d39;
		889: SAMPLE = 16'h7d43;
		890: SAMPLE = 16'h7d4e;
		891: SAMPLE = 16'h7d58;
		892: SAMPLE = 16'h7d62;
		893: SAMPLE = 16'h7d6c;
		894: SAMPLE = 16'h7d76;
		895: SAMPLE = 16'h7d80;
		896: SAMPLE = 16'h7d8a;
		897: SAMPLE = 16'h7d94;
		898: SAMPLE = 16'h7d9d;
		899: SAMPLE = 16'h7da7;
		900: SAMPLE = 16'h7db0;
		901: SAMPLE = 16'h7dba;
		902: SAMPLE = 16'h7dc3;
		903: SAMPLE = 16'h7dcd;
		904: SAMPLE = 16'h7dd6;
		905: SAMPLE = 16'h7ddf;
		906: SAMPLE = 16'h7de8;
		907: SAMPLE = 16'h7df1;
		908: SAMPLE = 16'h7dfa;
		909: SAMPLE = 16'h7e03;
		910: SAMPLE = 16'h7e0c;
		911: SAMPLE = 16'h7e14;
		912: SAMPLE = 16'h7e1d;
		913: SAMPLE = 16'h7e26;
		914: SAMPLE = 16'h7e2e;
		915: SAMPLE = 16'h7e37;
		916: SAMPLE = 16'h7e3f;
		917: SAMPLE = 16'h7e47;
		918: SAMPLE = 16'h7e4f;
		919: SAMPLE = 16'h7e57;
		920: SAMPLE = 16'h7e5f;
		921: SAMPLE = 16'h7e67;
		922: SAMPLE = 16'h7e6f;
		923: SAMPLE = 16'h7e77;
		924: SAMPLE = 16'h7e7f;
		925: SAMPLE = 16'h7e86;
		926: SAMPLE = 16'h7e8e;
		927: SAMPLE = 16'h7e95;
		928: SAMPLE = 16'h7e9d;
		929: SAMPLE = 16'h7ea4;
		930: SAMPLE = 16'h7eab;
		931: SAMPLE = 16'h7eb3;
		932: SAMPLE = 16'h7eba;
		933: SAMPLE = 16'h7ec1;
		934: SAMPLE = 16'h7ec8;
		935: SAMPLE = 16'h7ecf;
		936: SAMPLE = 16'h7ed5;
		937: SAMPLE = 16'h7edc;
		938: SAMPLE = 16'h7ee3;
		939: SAMPLE = 16'h7ee9;
		940: SAMPLE = 16'h7ef0;
		941: SAMPLE = 16'h7ef6;
		942: SAMPLE = 16'h7efd;
		943: SAMPLE = 16'h7f03;
		944: SAMPLE = 16'h7f09;
		945: SAMPLE = 16'h7f0f;
		946: SAMPLE = 16'h7f15;
		947: SAMPLE = 16'h7f1b;
		948: SAMPLE = 16'h7f21;
		949: SAMPLE = 16'h7f27;
		950: SAMPLE = 16'h7f2d;
		951: SAMPLE = 16'h7f32;
		952: SAMPLE = 16'h7f38;
		953: SAMPLE = 16'h7f3d;
		954: SAMPLE = 16'h7f43;
		955: SAMPLE = 16'h7f48;
		956: SAMPLE = 16'h7f4d;
		957: SAMPLE = 16'h7f53;
		958: SAMPLE = 16'h7f58;
		959: SAMPLE = 16'h7f5d;
		960: SAMPLE = 16'h7f62;
		961: SAMPLE = 16'h7f67;
		962: SAMPLE = 16'h7f6b;
		963: SAMPLE = 16'h7f70;
		964: SAMPLE = 16'h7f75;
		965: SAMPLE = 16'h7f79;
		966: SAMPLE = 16'h7f7e;
		967: SAMPLE = 16'h7f82;
		968: SAMPLE = 16'h7f87;
		969: SAMPLE = 16'h7f8b;
		970: SAMPLE = 16'h7f8f;
		971: SAMPLE = 16'h7f93;
		972: SAMPLE = 16'h7f97;
		973: SAMPLE = 16'h7f9b;
		974: SAMPLE = 16'h7f9f;
		975: SAMPLE = 16'h7fa3;
		976: SAMPLE = 16'h7fa7;
		977: SAMPLE = 16'h7faa;
		978: SAMPLE = 16'h7fae;
		979: SAMPLE = 16'h7fb1;
		980: SAMPLE = 16'h7fb5;
		981: SAMPLE = 16'h7fb8;
		982: SAMPLE = 16'h7fbc;
		983: SAMPLE = 16'h7fbf;
		984: SAMPLE = 16'h7fc2;
		985: SAMPLE = 16'h7fc5;
		986: SAMPLE = 16'h7fc8;
		987: SAMPLE = 16'h7fcb;
		988: SAMPLE = 16'h7fce;
		989: SAMPLE = 16'h7fd0;
		990: SAMPLE = 16'h7fd3;
		991: SAMPLE = 16'h7fd6;
		992: SAMPLE = 16'h7fd8;
		993: SAMPLE = 16'h7fda;
		994: SAMPLE = 16'h7fdd;
		995: SAMPLE = 16'h7fdf;
		996: SAMPLE = 16'h7fe1;
		997: SAMPLE = 16'h7fe3;
		998: SAMPLE = 16'h7fe5;
		999: SAMPLE = 16'h7fe7;
		1000: SAMPLE = 16'h7fe9;
		1001: SAMPLE = 16'h7feb;
		1002: SAMPLE = 16'h7fed;
		1003: SAMPLE = 16'h7fee;
		1004: SAMPLE = 16'h7ff0;
		1005: SAMPLE = 16'h7ff2;
		1006: SAMPLE = 16'h7ff3;
		1007: SAMPLE = 16'h7ff4;
		1008: SAMPLE = 16'h7ff6;
		1009: SAMPLE = 16'h7ff7;
		1010: SAMPLE = 16'h7ff8;
		1011: SAMPLE = 16'h7ff9;
		1012: SAMPLE = 16'h7ffa;
		1013: SAMPLE = 16'h7ffb;
		1014: SAMPLE = 16'h7ffc;
		1015: SAMPLE = 16'h7ffc;
		1016: SAMPLE = 16'h7ffd;
		1017: SAMPLE = 16'h7ffe;
		1018: SAMPLE = 16'h7ffe;
		1019: SAMPLE = 16'h7fff;
		1020: SAMPLE = 16'h7fff;
		1021: SAMPLE = 16'h7fff;
		1022: SAMPLE = 16'h7fff;
		1023: SAMPLE = 16'h7fff;
		1024: SAMPLE = 16'h8000;
		1025: SAMPLE = 16'h7fff;
		1026: SAMPLE = 16'h7fff;
		1027: SAMPLE = 16'h7fff;
		1028: SAMPLE = 16'h7fff;
		1029: SAMPLE = 16'h7fff;
		1030: SAMPLE = 16'h7ffe;
		1031: SAMPLE = 16'h7ffe;
		1032: SAMPLE = 16'h7ffd;
		1033: SAMPLE = 16'h7ffc;
		1034: SAMPLE = 16'h7ffc;
		1035: SAMPLE = 16'h7ffb;
		1036: SAMPLE = 16'h7ffa;
		1037: SAMPLE = 16'h7ff9;
		1038: SAMPLE = 16'h7ff8;
		1039: SAMPLE = 16'h7ff7;
		1040: SAMPLE = 16'h7ff6;
		1041: SAMPLE = 16'h7ff4;
		1042: SAMPLE = 16'h7ff3;
		1043: SAMPLE = 16'h7ff2;
		1044: SAMPLE = 16'h7ff0;
		1045: SAMPLE = 16'h7fee;
		1046: SAMPLE = 16'h7fed;
		1047: SAMPLE = 16'h7feb;
		1048: SAMPLE = 16'h7fe9;
		1049: SAMPLE = 16'h7fe7;
		1050: SAMPLE = 16'h7fe5;
		1051: SAMPLE = 16'h7fe3;
		1052: SAMPLE = 16'h7fe1;
		1053: SAMPLE = 16'h7fdf;
		1054: SAMPLE = 16'h7fdd;
		1055: SAMPLE = 16'h7fda;
		1056: SAMPLE = 16'h7fd8;
		1057: SAMPLE = 16'h7fd6;
		1058: SAMPLE = 16'h7fd3;
		1059: SAMPLE = 16'h7fd0;
		1060: SAMPLE = 16'h7fce;
		1061: SAMPLE = 16'h7fcb;
		1062: SAMPLE = 16'h7fc8;
		1063: SAMPLE = 16'h7fc5;
		1064: SAMPLE = 16'h7fc2;
		1065: SAMPLE = 16'h7fbf;
		1066: SAMPLE = 16'h7fbc;
		1067: SAMPLE = 16'h7fb8;
		1068: SAMPLE = 16'h7fb5;
		1069: SAMPLE = 16'h7fb1;
		1070: SAMPLE = 16'h7fae;
		1071: SAMPLE = 16'h7faa;
		1072: SAMPLE = 16'h7fa7;
		1073: SAMPLE = 16'h7fa3;
		1074: SAMPLE = 16'h7f9f;
		1075: SAMPLE = 16'h7f9b;
		1076: SAMPLE = 16'h7f97;
		1077: SAMPLE = 16'h7f93;
		1078: SAMPLE = 16'h7f8f;
		1079: SAMPLE = 16'h7f8b;
		1080: SAMPLE = 16'h7f87;
		1081: SAMPLE = 16'h7f82;
		1082: SAMPLE = 16'h7f7e;
		1083: SAMPLE = 16'h7f79;
		1084: SAMPLE = 16'h7f75;
		1085: SAMPLE = 16'h7f70;
		1086: SAMPLE = 16'h7f6b;
		1087: SAMPLE = 16'h7f67;
		1088: SAMPLE = 16'h7f62;
		1089: SAMPLE = 16'h7f5d;
		1090: SAMPLE = 16'h7f58;
		1091: SAMPLE = 16'h7f53;
		1092: SAMPLE = 16'h7f4d;
		1093: SAMPLE = 16'h7f48;
		1094: SAMPLE = 16'h7f43;
		1095: SAMPLE = 16'h7f3d;
		1096: SAMPLE = 16'h7f38;
		1097: SAMPLE = 16'h7f32;
		1098: SAMPLE = 16'h7f2d;
		1099: SAMPLE = 16'h7f27;
		1100: SAMPLE = 16'h7f21;
		1101: SAMPLE = 16'h7f1b;
		1102: SAMPLE = 16'h7f15;
		1103: SAMPLE = 16'h7f0f;
		1104: SAMPLE = 16'h7f09;
		1105: SAMPLE = 16'h7f03;
		1106: SAMPLE = 16'h7efd;
		1107: SAMPLE = 16'h7ef6;
		1108: SAMPLE = 16'h7ef0;
		1109: SAMPLE = 16'h7ee9;
		1110: SAMPLE = 16'h7ee3;
		1111: SAMPLE = 16'h7edc;
		1112: SAMPLE = 16'h7ed5;
		1113: SAMPLE = 16'h7ecf;
		1114: SAMPLE = 16'h7ec8;
		1115: SAMPLE = 16'h7ec1;
		1116: SAMPLE = 16'h7eba;
		1117: SAMPLE = 16'h7eb3;
		1118: SAMPLE = 16'h7eab;
		1119: SAMPLE = 16'h7ea4;
		1120: SAMPLE = 16'h7e9d;
		1121: SAMPLE = 16'h7e95;
		1122: SAMPLE = 16'h7e8e;
		1123: SAMPLE = 16'h7e86;
		1124: SAMPLE = 16'h7e7f;
		1125: SAMPLE = 16'h7e77;
		1126: SAMPLE = 16'h7e6f;
		1127: SAMPLE = 16'h7e67;
		1128: SAMPLE = 16'h7e5f;
		1129: SAMPLE = 16'h7e57;
		1130: SAMPLE = 16'h7e4f;
		1131: SAMPLE = 16'h7e47;
		1132: SAMPLE = 16'h7e3f;
		1133: SAMPLE = 16'h7e37;
		1134: SAMPLE = 16'h7e2e;
		1135: SAMPLE = 16'h7e26;
		1136: SAMPLE = 16'h7e1d;
		1137: SAMPLE = 16'h7e14;
		1138: SAMPLE = 16'h7e0c;
		1139: SAMPLE = 16'h7e03;
		1140: SAMPLE = 16'h7dfa;
		1141: SAMPLE = 16'h7df1;
		1142: SAMPLE = 16'h7de8;
		1143: SAMPLE = 16'h7ddf;
		1144: SAMPLE = 16'h7dd6;
		1145: SAMPLE = 16'h7dcd;
		1146: SAMPLE = 16'h7dc3;
		1147: SAMPLE = 16'h7dba;
		1148: SAMPLE = 16'h7db0;
		1149: SAMPLE = 16'h7da7;
		1150: SAMPLE = 16'h7d9d;
		1151: SAMPLE = 16'h7d94;
		1152: SAMPLE = 16'h7d8a;
		1153: SAMPLE = 16'h7d80;
		1154: SAMPLE = 16'h7d76;
		1155: SAMPLE = 16'h7d6c;
		1156: SAMPLE = 16'h7d62;
		1157: SAMPLE = 16'h7d58;
		1158: SAMPLE = 16'h7d4e;
		1159: SAMPLE = 16'h7d43;
		1160: SAMPLE = 16'h7d39;
		1161: SAMPLE = 16'h7d2f;
		1162: SAMPLE = 16'h7d24;
		1163: SAMPLE = 16'h7d19;
		1164: SAMPLE = 16'h7d0f;
		1165: SAMPLE = 16'h7d04;
		1166: SAMPLE = 16'h7cf9;
		1167: SAMPLE = 16'h7cee;
		1168: SAMPLE = 16'h7ce3;
		1169: SAMPLE = 16'h7cd8;
		1170: SAMPLE = 16'h7ccd;
		1171: SAMPLE = 16'h7cc2;
		1172: SAMPLE = 16'h7cb7;
		1173: SAMPLE = 16'h7cab;
		1174: SAMPLE = 16'h7ca0;
		1175: SAMPLE = 16'h7c94;
		1176: SAMPLE = 16'h7c89;
		1177: SAMPLE = 16'h7c7d;
		1178: SAMPLE = 16'h7c71;
		1179: SAMPLE = 16'h7c66;
		1180: SAMPLE = 16'h7c5a;
		1181: SAMPLE = 16'h7c4e;
		1182: SAMPLE = 16'h7c42;
		1183: SAMPLE = 16'h7c36;
		1184: SAMPLE = 16'h7c29;
		1185: SAMPLE = 16'h7c1d;
		1186: SAMPLE = 16'h7c11;
		1187: SAMPLE = 16'h7c05;
		1188: SAMPLE = 16'h7bf8;
		1189: SAMPLE = 16'h7beb;
		1190: SAMPLE = 16'h7bdf;
		1191: SAMPLE = 16'h7bd2;
		1192: SAMPLE = 16'h7bc5;
		1193: SAMPLE = 16'h7bb9;
		1194: SAMPLE = 16'h7bac;
		1195: SAMPLE = 16'h7b9f;
		1196: SAMPLE = 16'h7b92;
		1197: SAMPLE = 16'h7b84;
		1198: SAMPLE = 16'h7b77;
		1199: SAMPLE = 16'h7b6a;
		1200: SAMPLE = 16'h7b5d;
		1201: SAMPLE = 16'h7b4f;
		1202: SAMPLE = 16'h7b42;
		1203: SAMPLE = 16'h7b34;
		1204: SAMPLE = 16'h7b26;
		1205: SAMPLE = 16'h7b19;
		1206: SAMPLE = 16'h7b0b;
		1207: SAMPLE = 16'h7afd;
		1208: SAMPLE = 16'h7aef;
		1209: SAMPLE = 16'h7ae1;
		1210: SAMPLE = 16'h7ad3;
		1211: SAMPLE = 16'h7ac5;
		1212: SAMPLE = 16'h7ab6;
		1213: SAMPLE = 16'h7aa8;
		1214: SAMPLE = 16'h7a9a;
		1215: SAMPLE = 16'h7a8b;
		1216: SAMPLE = 16'h7a7d;
		1217: SAMPLE = 16'h7a6e;
		1218: SAMPLE = 16'h7a5f;
		1219: SAMPLE = 16'h7a50;
		1220: SAMPLE = 16'h7a42;
		1221: SAMPLE = 16'h7a33;
		1222: SAMPLE = 16'h7a24;
		1223: SAMPLE = 16'h7a15;
		1224: SAMPLE = 16'h7a05;
		1225: SAMPLE = 16'h79f6;
		1226: SAMPLE = 16'h79e7;
		1227: SAMPLE = 16'h79d8;
		1228: SAMPLE = 16'h79c8;
		1229: SAMPLE = 16'h79b9;
		1230: SAMPLE = 16'h79a9;
		1231: SAMPLE = 16'h7999;
		1232: SAMPLE = 16'h798a;
		1233: SAMPLE = 16'h797a;
		1234: SAMPLE = 16'h796a;
		1235: SAMPLE = 16'h795a;
		1236: SAMPLE = 16'h794a;
		1237: SAMPLE = 16'h793a;
		1238: SAMPLE = 16'h792a;
		1239: SAMPLE = 16'h7919;
		1240: SAMPLE = 16'h7909;
		1241: SAMPLE = 16'h78f9;
		1242: SAMPLE = 16'h78e8;
		1243: SAMPLE = 16'h78d8;
		1244: SAMPLE = 16'h78c7;
		1245: SAMPLE = 16'h78b6;
		1246: SAMPLE = 16'h78a6;
		1247: SAMPLE = 16'h7895;
		1248: SAMPLE = 16'h7884;
		1249: SAMPLE = 16'h7873;
		1250: SAMPLE = 16'h7862;
		1251: SAMPLE = 16'h7851;
		1252: SAMPLE = 16'h7840;
		1253: SAMPLE = 16'h782e;
		1254: SAMPLE = 16'h781d;
		1255: SAMPLE = 16'h780c;
		1256: SAMPLE = 16'h77fa;
		1257: SAMPLE = 16'h77e9;
		1258: SAMPLE = 16'h77d7;
		1259: SAMPLE = 16'h77c5;
		1260: SAMPLE = 16'h77b4;
		1261: SAMPLE = 16'h77a2;
		1262: SAMPLE = 16'h7790;
		1263: SAMPLE = 16'h777e;
		1264: SAMPLE = 16'h776c;
		1265: SAMPLE = 16'h775a;
		1266: SAMPLE = 16'h7747;
		1267: SAMPLE = 16'h7735;
		1268: SAMPLE = 16'h7723;
		1269: SAMPLE = 16'h7710;
		1270: SAMPLE = 16'h76fe;
		1271: SAMPLE = 16'h76eb;
		1272: SAMPLE = 16'h76d9;
		1273: SAMPLE = 16'h76c6;
		1274: SAMPLE = 16'h76b3;
		1275: SAMPLE = 16'h76a0;
		1276: SAMPLE = 16'h768e;
		1277: SAMPLE = 16'h767b;
		1278: SAMPLE = 16'h7668;
		1279: SAMPLE = 16'h7654;
		1280: SAMPLE = 16'h7641;
		1281: SAMPLE = 16'h762e;
		1282: SAMPLE = 16'h761b;
		1283: SAMPLE = 16'h7607;
		1284: SAMPLE = 16'h75f4;
		1285: SAMPLE = 16'h75e0;
		1286: SAMPLE = 16'h75cc;
		1287: SAMPLE = 16'h75b9;
		1288: SAMPLE = 16'h75a5;
		1289: SAMPLE = 16'h7591;
		1290: SAMPLE = 16'h757d;
		1291: SAMPLE = 16'h7569;
		1292: SAMPLE = 16'h7555;
		1293: SAMPLE = 16'h7541;
		1294: SAMPLE = 16'h752d;
		1295: SAMPLE = 16'h7519;
		1296: SAMPLE = 16'h7504;
		1297: SAMPLE = 16'h74f0;
		1298: SAMPLE = 16'h74db;
		1299: SAMPLE = 16'h74c7;
		1300: SAMPLE = 16'h74b2;
		1301: SAMPLE = 16'h749e;
		1302: SAMPLE = 16'h7489;
		1303: SAMPLE = 16'h7474;
		1304: SAMPLE = 16'h745f;
		1305: SAMPLE = 16'h744a;
		1306: SAMPLE = 16'h7435;
		1307: SAMPLE = 16'h7420;
		1308: SAMPLE = 16'h740b;
		1309: SAMPLE = 16'h73f6;
		1310: SAMPLE = 16'h73e0;
		1311: SAMPLE = 16'h73cb;
		1312: SAMPLE = 16'h73b5;
		1313: SAMPLE = 16'h73a0;
		1314: SAMPLE = 16'h738a;
		1315: SAMPLE = 16'h7375;
		1316: SAMPLE = 16'h735f;
		1317: SAMPLE = 16'h7349;
		1318: SAMPLE = 16'h7333;
		1319: SAMPLE = 16'h731d;
		1320: SAMPLE = 16'h7307;
		1321: SAMPLE = 16'h72f1;
		1322: SAMPLE = 16'h72db;
		1323: SAMPLE = 16'h72c5;
		1324: SAMPLE = 16'h72af;
		1325: SAMPLE = 16'h7298;
		1326: SAMPLE = 16'h7282;
		1327: SAMPLE = 16'h726b;
		1328: SAMPLE = 16'h7255;
		1329: SAMPLE = 16'h723e;
		1330: SAMPLE = 16'h7227;
		1331: SAMPLE = 16'h7211;
		1332: SAMPLE = 16'h71fa;
		1333: SAMPLE = 16'h71e3;
		1334: SAMPLE = 16'h71cc;
		1335: SAMPLE = 16'h71b5;
		1336: SAMPLE = 16'h719e;
		1337: SAMPLE = 16'h7186;
		1338: SAMPLE = 16'h716f;
		1339: SAMPLE = 16'h7158;
		1340: SAMPLE = 16'h7141;
		1341: SAMPLE = 16'h7129;
		1342: SAMPLE = 16'h7112;
		1343: SAMPLE = 16'h70fa;
		1344: SAMPLE = 16'h70e2;
		1345: SAMPLE = 16'h70cb;
		1346: SAMPLE = 16'h70b3;
		1347: SAMPLE = 16'h709b;
		1348: SAMPLE = 16'h7083;
		1349: SAMPLE = 16'h706b;
		1350: SAMPLE = 16'h7053;
		1351: SAMPLE = 16'h703b;
		1352: SAMPLE = 16'h7023;
		1353: SAMPLE = 16'h700a;
		1354: SAMPLE = 16'h6ff2;
		1355: SAMPLE = 16'h6fda;
		1356: SAMPLE = 16'h6fc1;
		1357: SAMPLE = 16'h6fa9;
		1358: SAMPLE = 16'h6f90;
		1359: SAMPLE = 16'h6f77;
		1360: SAMPLE = 16'h6f5f;
		1361: SAMPLE = 16'h6f46;
		1362: SAMPLE = 16'h6f2d;
		1363: SAMPLE = 16'h6f14;
		1364: SAMPLE = 16'h6efb;
		1365: SAMPLE = 16'h6ee2;
		1366: SAMPLE = 16'h6ec9;
		1367: SAMPLE = 16'h6eaf;
		1368: SAMPLE = 16'h6e96;
		1369: SAMPLE = 16'h6e7d;
		1370: SAMPLE = 16'h6e63;
		1371: SAMPLE = 16'h6e4a;
		1372: SAMPLE = 16'h6e30;
		1373: SAMPLE = 16'h6e17;
		1374: SAMPLE = 16'h6dfd;
		1375: SAMPLE = 16'h6de3;
		1376: SAMPLE = 16'h6dca;
		1377: SAMPLE = 16'h6db0;
		1378: SAMPLE = 16'h6d96;
		1379: SAMPLE = 16'h6d7c;
		1380: SAMPLE = 16'h6d62;
		1381: SAMPLE = 16'h6d48;
		1382: SAMPLE = 16'h6d2d;
		1383: SAMPLE = 16'h6d13;
		1384: SAMPLE = 16'h6cf9;
		1385: SAMPLE = 16'h6cde;
		1386: SAMPLE = 16'h6cc4;
		1387: SAMPLE = 16'h6ca9;
		1388: SAMPLE = 16'h6c8f;
		1389: SAMPLE = 16'h6c74;
		1390: SAMPLE = 16'h6c59;
		1391: SAMPLE = 16'h6c3f;
		1392: SAMPLE = 16'h6c24;
		1393: SAMPLE = 16'h6c09;
		1394: SAMPLE = 16'h6bee;
		1395: SAMPLE = 16'h6bd3;
		1396: SAMPLE = 16'h6bb8;
		1397: SAMPLE = 16'h6b9c;
		1398: SAMPLE = 16'h6b81;
		1399: SAMPLE = 16'h6b66;
		1400: SAMPLE = 16'h6b4a;
		1401: SAMPLE = 16'h6b2f;
		1402: SAMPLE = 16'h6b13;
		1403: SAMPLE = 16'h6af8;
		1404: SAMPLE = 16'h6adc;
		1405: SAMPLE = 16'h6ac1;
		1406: SAMPLE = 16'h6aa5;
		1407: SAMPLE = 16'h6a89;
		1408: SAMPLE = 16'h6a6d;
		1409: SAMPLE = 16'h6a51;
		1410: SAMPLE = 16'h6a35;
		1411: SAMPLE = 16'h6a19;
		1412: SAMPLE = 16'h69fd;
		1413: SAMPLE = 16'h69e1;
		1414: SAMPLE = 16'h69c4;
		1415: SAMPLE = 16'h69a8;
		1416: SAMPLE = 16'h698c;
		1417: SAMPLE = 16'h696f;
		1418: SAMPLE = 16'h6953;
		1419: SAMPLE = 16'h6936;
		1420: SAMPLE = 16'h6919;
		1421: SAMPLE = 16'h68fd;
		1422: SAMPLE = 16'h68e0;
		1423: SAMPLE = 16'h68c3;
		1424: SAMPLE = 16'h68a6;
		1425: SAMPLE = 16'h6889;
		1426: SAMPLE = 16'h686c;
		1427: SAMPLE = 16'h684f;
		1428: SAMPLE = 16'h6832;
		1429: SAMPLE = 16'h6815;
		1430: SAMPLE = 16'h67f7;
		1431: SAMPLE = 16'h67da;
		1432: SAMPLE = 16'h67bd;
		1433: SAMPLE = 16'h679f;
		1434: SAMPLE = 16'h6782;
		1435: SAMPLE = 16'h6764;
		1436: SAMPLE = 16'h6746;
		1437: SAMPLE = 16'h6729;
		1438: SAMPLE = 16'h670b;
		1439: SAMPLE = 16'h66ed;
		1440: SAMPLE = 16'h66cf;
		1441: SAMPLE = 16'h66b1;
		1442: SAMPLE = 16'h6693;
		1443: SAMPLE = 16'h6675;
		1444: SAMPLE = 16'h6657;
		1445: SAMPLE = 16'h6639;
		1446: SAMPLE = 16'h661a;
		1447: SAMPLE = 16'h65fc;
		1448: SAMPLE = 16'h65dd;
		1449: SAMPLE = 16'h65bf;
		1450: SAMPLE = 16'h65a0;
		1451: SAMPLE = 16'h6582;
		1452: SAMPLE = 16'h6563;
		1453: SAMPLE = 16'h6545;
		1454: SAMPLE = 16'h6526;
		1455: SAMPLE = 16'h6507;
		1456: SAMPLE = 16'h64e8;
		1457: SAMPLE = 16'h64c9;
		1458: SAMPLE = 16'h64aa;
		1459: SAMPLE = 16'h648b;
		1460: SAMPLE = 16'h646c;
		1461: SAMPLE = 16'h644d;
		1462: SAMPLE = 16'h642d;
		1463: SAMPLE = 16'h640e;
		1464: SAMPLE = 16'h63ef;
		1465: SAMPLE = 16'h63cf;
		1466: SAMPLE = 16'h63b0;
		1467: SAMPLE = 16'h6390;
		1468: SAMPLE = 16'h6371;
		1469: SAMPLE = 16'h6351;
		1470: SAMPLE = 16'h6331;
		1471: SAMPLE = 16'h6311;
		1472: SAMPLE = 16'h62f2;
		1473: SAMPLE = 16'h62d2;
		1474: SAMPLE = 16'h62b2;
		1475: SAMPLE = 16'h6292;
		1476: SAMPLE = 16'h6271;
		1477: SAMPLE = 16'h6251;
		1478: SAMPLE = 16'h6231;
		1479: SAMPLE = 16'h6211;
		1480: SAMPLE = 16'h61f1;
		1481: SAMPLE = 16'h61d0;
		1482: SAMPLE = 16'h61b0;
		1483: SAMPLE = 16'h618f;
		1484: SAMPLE = 16'h616f;
		1485: SAMPLE = 16'h614e;
		1486: SAMPLE = 16'h612d;
		1487: SAMPLE = 16'h610d;
		1488: SAMPLE = 16'h60ec;
		1489: SAMPLE = 16'h60cb;
		1490: SAMPLE = 16'h60aa;
		1491: SAMPLE = 16'h6089;
		1492: SAMPLE = 16'h6068;
		1493: SAMPLE = 16'h6047;
		1494: SAMPLE = 16'h6026;
		1495: SAMPLE = 16'h6004;
		1496: SAMPLE = 16'h5fe3;
		1497: SAMPLE = 16'h5fc2;
		1498: SAMPLE = 16'h5fa0;
		1499: SAMPLE = 16'h5f7f;
		1500: SAMPLE = 16'h5f5e;
		1501: SAMPLE = 16'h5f3c;
		1502: SAMPLE = 16'h5f1a;
		1503: SAMPLE = 16'h5ef9;
		1504: SAMPLE = 16'h5ed7;
		1505: SAMPLE = 16'h5eb5;
		1506: SAMPLE = 16'h5e93;
		1507: SAMPLE = 16'h5e71;
		1508: SAMPLE = 16'h5e50;
		1509: SAMPLE = 16'h5e2d;
		1510: SAMPLE = 16'h5e0b;
		1511: SAMPLE = 16'h5de9;
		1512: SAMPLE = 16'h5dc7;
		1513: SAMPLE = 16'h5da5;
		1514: SAMPLE = 16'h5d83;
		1515: SAMPLE = 16'h5d60;
		1516: SAMPLE = 16'h5d3e;
		1517: SAMPLE = 16'h5d1b;
		1518: SAMPLE = 16'h5cf9;
		1519: SAMPLE = 16'h5cd6;
		1520: SAMPLE = 16'h5cb4;
		1521: SAMPLE = 16'h5c91;
		1522: SAMPLE = 16'h5c6e;
		1523: SAMPLE = 16'h5c4b;
		1524: SAMPLE = 16'h5c29;
		1525: SAMPLE = 16'h5c06;
		1526: SAMPLE = 16'h5be3;
		1527: SAMPLE = 16'h5bc0;
		1528: SAMPLE = 16'h5b9d;
		1529: SAMPLE = 16'h5b79;
		1530: SAMPLE = 16'h5b56;
		1531: SAMPLE = 16'h5b33;
		1532: SAMPLE = 16'h5b10;
		1533: SAMPLE = 16'h5aec;
		1534: SAMPLE = 16'h5ac9;
		1535: SAMPLE = 16'h5aa5;
		1536: SAMPLE = 16'h5a82;
		1537: SAMPLE = 16'h5a5e;
		1538: SAMPLE = 16'h5a3b;
		1539: SAMPLE = 16'h5a17;
		1540: SAMPLE = 16'h59f3;
		1541: SAMPLE = 16'h59d0;
		1542: SAMPLE = 16'h59ac;
		1543: SAMPLE = 16'h5988;
		1544: SAMPLE = 16'h5964;
		1545: SAMPLE = 16'h5940;
		1546: SAMPLE = 16'h591c;
		1547: SAMPLE = 16'h58f8;
		1548: SAMPLE = 16'h58d4;
		1549: SAMPLE = 16'h58af;
		1550: SAMPLE = 16'h588b;
		1551: SAMPLE = 16'h5867;
		1552: SAMPLE = 16'h5842;
		1553: SAMPLE = 16'h581e;
		1554: SAMPLE = 16'h57f9;
		1555: SAMPLE = 16'h57d5;
		1556: SAMPLE = 16'h57b0;
		1557: SAMPLE = 16'h578c;
		1558: SAMPLE = 16'h5767;
		1559: SAMPLE = 16'h5742;
		1560: SAMPLE = 16'h571d;
		1561: SAMPLE = 16'h56f9;
		1562: SAMPLE = 16'h56d4;
		1563: SAMPLE = 16'h56af;
		1564: SAMPLE = 16'h568a;
		1565: SAMPLE = 16'h5665;
		1566: SAMPLE = 16'h5640;
		1567: SAMPLE = 16'h561a;
		1568: SAMPLE = 16'h55f5;
		1569: SAMPLE = 16'h55d0;
		1570: SAMPLE = 16'h55ab;
		1571: SAMPLE = 16'h5585;
		1572: SAMPLE = 16'h5560;
		1573: SAMPLE = 16'h553a;
		1574: SAMPLE = 16'h5515;
		1575: SAMPLE = 16'h54ef;
		1576: SAMPLE = 16'h54ca;
		1577: SAMPLE = 16'h54a4;
		1578: SAMPLE = 16'h547e;
		1579: SAMPLE = 16'h5458;
		1580: SAMPLE = 16'h5433;
		1581: SAMPLE = 16'h540d;
		1582: SAMPLE = 16'h53e7;
		1583: SAMPLE = 16'h53c1;
		1584: SAMPLE = 16'h539b;
		1585: SAMPLE = 16'h5375;
		1586: SAMPLE = 16'h534e;
		1587: SAMPLE = 16'h5328;
		1588: SAMPLE = 16'h5302;
		1589: SAMPLE = 16'h52dc;
		1590: SAMPLE = 16'h52b5;
		1591: SAMPLE = 16'h528f;
		1592: SAMPLE = 16'h5269;
		1593: SAMPLE = 16'h5242;
		1594: SAMPLE = 16'h521c;
		1595: SAMPLE = 16'h51f5;
		1596: SAMPLE = 16'h51ce;
		1597: SAMPLE = 16'h51a8;
		1598: SAMPLE = 16'h5181;
		1599: SAMPLE = 16'h515a;
		1600: SAMPLE = 16'h5133;
		1601: SAMPLE = 16'h510c;
		1602: SAMPLE = 16'h50e5;
		1603: SAMPLE = 16'h50bf;
		1604: SAMPLE = 16'h5097;
		1605: SAMPLE = 16'h5070;
		1606: SAMPLE = 16'h5049;
		1607: SAMPLE = 16'h5022;
		1608: SAMPLE = 16'h4ffb;
		1609: SAMPLE = 16'h4fd4;
		1610: SAMPLE = 16'h4fac;
		1611: SAMPLE = 16'h4f85;
		1612: SAMPLE = 16'h4f5e;
		1613: SAMPLE = 16'h4f36;
		1614: SAMPLE = 16'h4f0f;
		1615: SAMPLE = 16'h4ee7;
		1616: SAMPLE = 16'h4ebf;
		1617: SAMPLE = 16'h4e98;
		1618: SAMPLE = 16'h4e70;
		1619: SAMPLE = 16'h4e48;
		1620: SAMPLE = 16'h4e21;
		1621: SAMPLE = 16'h4df9;
		1622: SAMPLE = 16'h4dd1;
		1623: SAMPLE = 16'h4da9;
		1624: SAMPLE = 16'h4d81;
		1625: SAMPLE = 16'h4d59;
		1626: SAMPLE = 16'h4d31;
		1627: SAMPLE = 16'h4d09;
		1628: SAMPLE = 16'h4ce1;
		1629: SAMPLE = 16'h4cb8;
		1630: SAMPLE = 16'h4c90;
		1631: SAMPLE = 16'h4c68;
		1632: SAMPLE = 16'h4c3f;
		1633: SAMPLE = 16'h4c17;
		1634: SAMPLE = 16'h4bef;
		1635: SAMPLE = 16'h4bc6;
		1636: SAMPLE = 16'h4b9e;
		1637: SAMPLE = 16'h4b75;
		1638: SAMPLE = 16'h4b4c;
		1639: SAMPLE = 16'h4b24;
		1640: SAMPLE = 16'h4afb;
		1641: SAMPLE = 16'h4ad2;
		1642: SAMPLE = 16'h4aa9;
		1643: SAMPLE = 16'h4a81;
		1644: SAMPLE = 16'h4a58;
		1645: SAMPLE = 16'h4a2f;
		1646: SAMPLE = 16'h4a06;
		1647: SAMPLE = 16'h49dd;
		1648: SAMPLE = 16'h49b4;
		1649: SAMPLE = 16'h498a;
		1650: SAMPLE = 16'h4961;
		1651: SAMPLE = 16'h4938;
		1652: SAMPLE = 16'h490f;
		1653: SAMPLE = 16'h48e6;
		1654: SAMPLE = 16'h48bc;
		1655: SAMPLE = 16'h4893;
		1656: SAMPLE = 16'h4869;
		1657: SAMPLE = 16'h4840;
		1658: SAMPLE = 16'h4816;
		1659: SAMPLE = 16'h47ed;
		1660: SAMPLE = 16'h47c3;
		1661: SAMPLE = 16'h479a;
		1662: SAMPLE = 16'h4770;
		1663: SAMPLE = 16'h4746;
		1664: SAMPLE = 16'h471c;
		1665: SAMPLE = 16'h46f3;
		1666: SAMPLE = 16'h46c9;
		1667: SAMPLE = 16'h469f;
		1668: SAMPLE = 16'h4675;
		1669: SAMPLE = 16'h464b;
		1670: SAMPLE = 16'h4621;
		1671: SAMPLE = 16'h45f7;
		1672: SAMPLE = 16'h45cd;
		1673: SAMPLE = 16'h45a3;
		1674: SAMPLE = 16'h4578;
		1675: SAMPLE = 16'h454e;
		1676: SAMPLE = 16'h4524;
		1677: SAMPLE = 16'h44fa;
		1678: SAMPLE = 16'h44cf;
		1679: SAMPLE = 16'h44a5;
		1680: SAMPLE = 16'h447a;
		1681: SAMPLE = 16'h4450;
		1682: SAMPLE = 16'h4425;
		1683: SAMPLE = 16'h43fb;
		1684: SAMPLE = 16'h43d0;
		1685: SAMPLE = 16'h43a5;
		1686: SAMPLE = 16'h437b;
		1687: SAMPLE = 16'h4350;
		1688: SAMPLE = 16'h4325;
		1689: SAMPLE = 16'h42fa;
		1690: SAMPLE = 16'h42d0;
		1691: SAMPLE = 16'h42a5;
		1692: SAMPLE = 16'h427a;
		1693: SAMPLE = 16'h424f;
		1694: SAMPLE = 16'h4224;
		1695: SAMPLE = 16'h41f9;
		1696: SAMPLE = 16'h41ce;
		1697: SAMPLE = 16'h41a2;
		1698: SAMPLE = 16'h4177;
		1699: SAMPLE = 16'h414c;
		1700: SAMPLE = 16'h4121;
		1701: SAMPLE = 16'h40f6;
		1702: SAMPLE = 16'h40ca;
		1703: SAMPLE = 16'h409f;
		1704: SAMPLE = 16'h4073;
		1705: SAMPLE = 16'h4048;
		1706: SAMPLE = 16'h401d;
		1707: SAMPLE = 16'h3ff1;
		1708: SAMPLE = 16'h3fc5;
		1709: SAMPLE = 16'h3f9a;
		1710: SAMPLE = 16'h3f6e;
		1711: SAMPLE = 16'h3f43;
		1712: SAMPLE = 16'h3f17;
		1713: SAMPLE = 16'h3eeb;
		1714: SAMPLE = 16'h3ebf;
		1715: SAMPLE = 16'h3e93;
		1716: SAMPLE = 16'h3e68;
		1717: SAMPLE = 16'h3e3c;
		1718: SAMPLE = 16'h3e10;
		1719: SAMPLE = 16'h3de4;
		1720: SAMPLE = 16'h3db8;
		1721: SAMPLE = 16'h3d8c;
		1722: SAMPLE = 16'h3d60;
		1723: SAMPLE = 16'h3d33;
		1724: SAMPLE = 16'h3d07;
		1725: SAMPLE = 16'h3cdb;
		1726: SAMPLE = 16'h3caf;
		1727: SAMPLE = 16'h3c83;
		1728: SAMPLE = 16'h3c56;
		1729: SAMPLE = 16'h3c2a;
		1730: SAMPLE = 16'h3bfd;
		1731: SAMPLE = 16'h3bd1;
		1732: SAMPLE = 16'h3ba5;
		1733: SAMPLE = 16'h3b78;
		1734: SAMPLE = 16'h3b4c;
		1735: SAMPLE = 16'h3b1f;
		1736: SAMPLE = 16'h3af2;
		1737: SAMPLE = 16'h3ac6;
		1738: SAMPLE = 16'h3a99;
		1739: SAMPLE = 16'h3a6c;
		1740: SAMPLE = 16'h3a40;
		1741: SAMPLE = 16'h3a13;
		1742: SAMPLE = 16'h39e6;
		1743: SAMPLE = 16'h39b9;
		1744: SAMPLE = 16'h398c;
		1745: SAMPLE = 16'h395f;
		1746: SAMPLE = 16'h3932;
		1747: SAMPLE = 16'h3906;
		1748: SAMPLE = 16'h38d8;
		1749: SAMPLE = 16'h38ab;
		1750: SAMPLE = 16'h387e;
		1751: SAMPLE = 16'h3851;
		1752: SAMPLE = 16'h3824;
		1753: SAMPLE = 16'h37f7;
		1754: SAMPLE = 16'h37ca;
		1755: SAMPLE = 16'h379c;
		1756: SAMPLE = 16'h376f;
		1757: SAMPLE = 16'h3742;
		1758: SAMPLE = 16'h3714;
		1759: SAMPLE = 16'h36e7;
		1760: SAMPLE = 16'h36ba;
		1761: SAMPLE = 16'h368c;
		1762: SAMPLE = 16'h365f;
		1763: SAMPLE = 16'h3631;
		1764: SAMPLE = 16'h3604;
		1765: SAMPLE = 16'h35d6;
		1766: SAMPLE = 16'h35a8;
		1767: SAMPLE = 16'h357b;
		1768: SAMPLE = 16'h354d;
		1769: SAMPLE = 16'h351f;
		1770: SAMPLE = 16'h34f2;
		1771: SAMPLE = 16'h34c4;
		1772: SAMPLE = 16'h3496;
		1773: SAMPLE = 16'h3468;
		1774: SAMPLE = 16'h343a;
		1775: SAMPLE = 16'h340c;
		1776: SAMPLE = 16'h33de;
		1777: SAMPLE = 16'h33b0;
		1778: SAMPLE = 16'h3382;
		1779: SAMPLE = 16'h3354;
		1780: SAMPLE = 16'h3326;
		1781: SAMPLE = 16'h32f8;
		1782: SAMPLE = 16'h32ca;
		1783: SAMPLE = 16'h329c;
		1784: SAMPLE = 16'h326e;
		1785: SAMPLE = 16'h3240;
		1786: SAMPLE = 16'h3211;
		1787: SAMPLE = 16'h31e3;
		1788: SAMPLE = 16'h31b5;
		1789: SAMPLE = 16'h3186;
		1790: SAMPLE = 16'h3158;
		1791: SAMPLE = 16'h312a;
		1792: SAMPLE = 16'h30fb;
		1793: SAMPLE = 16'h30cd;
		1794: SAMPLE = 16'h309e;
		1795: SAMPLE = 16'h3070;
		1796: SAMPLE = 16'h3041;
		1797: SAMPLE = 16'h3013;
		1798: SAMPLE = 16'h2fe4;
		1799: SAMPLE = 16'h2fb5;
		1800: SAMPLE = 16'h2f87;
		1801: SAMPLE = 16'h2f58;
		1802: SAMPLE = 16'h2f29;
		1803: SAMPLE = 16'h2efb;
		1804: SAMPLE = 16'h2ecc;
		1805: SAMPLE = 16'h2e9d;
		1806: SAMPLE = 16'h2e6e;
		1807: SAMPLE = 16'h2e3f;
		1808: SAMPLE = 16'h2e11;
		1809: SAMPLE = 16'h2de2;
		1810: SAMPLE = 16'h2db3;
		1811: SAMPLE = 16'h2d84;
		1812: SAMPLE = 16'h2d55;
		1813: SAMPLE = 16'h2d26;
		1814: SAMPLE = 16'h2cf7;
		1815: SAMPLE = 16'h2cc8;
		1816: SAMPLE = 16'h2c98;
		1817: SAMPLE = 16'h2c69;
		1818: SAMPLE = 16'h2c3a;
		1819: SAMPLE = 16'h2c0b;
		1820: SAMPLE = 16'h2bdc;
		1821: SAMPLE = 16'h2bad;
		1822: SAMPLE = 16'h2b7d;
		1823: SAMPLE = 16'h2b4e;
		1824: SAMPLE = 16'h2b1f;
		1825: SAMPLE = 16'h2aef;
		1826: SAMPLE = 16'h2ac0;
		1827: SAMPLE = 16'h2a91;
		1828: SAMPLE = 16'h2a61;
		1829: SAMPLE = 16'h2a32;
		1830: SAMPLE = 16'h2a02;
		1831: SAMPLE = 16'h29d3;
		1832: SAMPLE = 16'h29a3;
		1833: SAMPLE = 16'h2974;
		1834: SAMPLE = 16'h2944;
		1835: SAMPLE = 16'h2915;
		1836: SAMPLE = 16'h28e5;
		1837: SAMPLE = 16'h28b5;
		1838: SAMPLE = 16'h2886;
		1839: SAMPLE = 16'h2856;
		1840: SAMPLE = 16'h2826;
		1841: SAMPLE = 16'h27f6;
		1842: SAMPLE = 16'h27c7;
		1843: SAMPLE = 16'h2797;
		1844: SAMPLE = 16'h2767;
		1845: SAMPLE = 16'h2737;
		1846: SAMPLE = 16'h2707;
		1847: SAMPLE = 16'h26d8;
		1848: SAMPLE = 16'h26a8;
		1849: SAMPLE = 16'h2678;
		1850: SAMPLE = 16'h2648;
		1851: SAMPLE = 16'h2618;
		1852: SAMPLE = 16'h25e8;
		1853: SAMPLE = 16'h25b8;
		1854: SAMPLE = 16'h2588;
		1855: SAMPLE = 16'h2558;
		1856: SAMPLE = 16'h2528;
		1857: SAMPLE = 16'h24f7;
		1858: SAMPLE = 16'h24c7;
		1859: SAMPLE = 16'h2497;
		1860: SAMPLE = 16'h2467;
		1861: SAMPLE = 16'h2437;
		1862: SAMPLE = 16'h2407;
		1863: SAMPLE = 16'h23d6;
		1864: SAMPLE = 16'h23a6;
		1865: SAMPLE = 16'h2376;
		1866: SAMPLE = 16'h2345;
		1867: SAMPLE = 16'h2315;
		1868: SAMPLE = 16'h22e5;
		1869: SAMPLE = 16'h22b4;
		1870: SAMPLE = 16'h2284;
		1871: SAMPLE = 16'h2254;
		1872: SAMPLE = 16'h2223;
		1873: SAMPLE = 16'h21f3;
		1874: SAMPLE = 16'h21c2;
		1875: SAMPLE = 16'h2192;
		1876: SAMPLE = 16'h2161;
		1877: SAMPLE = 16'h2131;
		1878: SAMPLE = 16'h2100;
		1879: SAMPLE = 16'h20d0;
		1880: SAMPLE = 16'h209f;
		1881: SAMPLE = 16'h206e;
		1882: SAMPLE = 16'h203e;
		1883: SAMPLE = 16'h200d;
		1884: SAMPLE = 16'h1fdc;
		1885: SAMPLE = 16'h1fac;
		1886: SAMPLE = 16'h1f7b;
		1887: SAMPLE = 16'h1f4a;
		1888: SAMPLE = 16'h1f19;
		1889: SAMPLE = 16'h1ee9;
		1890: SAMPLE = 16'h1eb8;
		1891: SAMPLE = 16'h1e87;
		1892: SAMPLE = 16'h1e56;
		1893: SAMPLE = 16'h1e25;
		1894: SAMPLE = 16'h1df5;
		1895: SAMPLE = 16'h1dc4;
		1896: SAMPLE = 16'h1d93;
		1897: SAMPLE = 16'h1d62;
		1898: SAMPLE = 16'h1d31;
		1899: SAMPLE = 16'h1d00;
		1900: SAMPLE = 16'h1ccf;
		1901: SAMPLE = 16'h1c9e;
		1902: SAMPLE = 16'h1c6d;
		1903: SAMPLE = 16'h1c3c;
		1904: SAMPLE = 16'h1c0b;
		1905: SAMPLE = 16'h1bda;
		1906: SAMPLE = 16'h1ba9;
		1907: SAMPLE = 16'h1b78;
		1908: SAMPLE = 16'h1b47;
		1909: SAMPLE = 16'h1b16;
		1910: SAMPLE = 16'h1ae4;
		1911: SAMPLE = 16'h1ab3;
		1912: SAMPLE = 16'h1a82;
		1913: SAMPLE = 16'h1a51;
		1914: SAMPLE = 16'h1a20;
		1915: SAMPLE = 16'h19ef;
		1916: SAMPLE = 16'h19bd;
		1917: SAMPLE = 16'h198c;
		1918: SAMPLE = 16'h195b;
		1919: SAMPLE = 16'h192a;
		1920: SAMPLE = 16'h18f8;
		1921: SAMPLE = 16'h18c7;
		1922: SAMPLE = 16'h1896;
		1923: SAMPLE = 16'h1864;
		1924: SAMPLE = 16'h1833;
		1925: SAMPLE = 16'h1802;
		1926: SAMPLE = 16'h17d0;
		1927: SAMPLE = 16'h179f;
		1928: SAMPLE = 16'h176d;
		1929: SAMPLE = 16'h173c;
		1930: SAMPLE = 16'h170a;
		1931: SAMPLE = 16'h16d9;
		1932: SAMPLE = 16'h16a8;
		1933: SAMPLE = 16'h1676;
		1934: SAMPLE = 16'h1645;
		1935: SAMPLE = 16'h1613;
		1936: SAMPLE = 16'h15e2;
		1937: SAMPLE = 16'h15b0;
		1938: SAMPLE = 16'h157f;
		1939: SAMPLE = 16'h154d;
		1940: SAMPLE = 16'h151b;
		1941: SAMPLE = 16'h14ea;
		1942: SAMPLE = 16'h14b8;
		1943: SAMPLE = 16'h1487;
		1944: SAMPLE = 16'h1455;
		1945: SAMPLE = 16'h1423;
		1946: SAMPLE = 16'h13f2;
		1947: SAMPLE = 16'h13c0;
		1948: SAMPLE = 16'h138e;
		1949: SAMPLE = 16'h135d;
		1950: SAMPLE = 16'h132b;
		1951: SAMPLE = 16'h12f9;
		1952: SAMPLE = 16'h12c8;
		1953: SAMPLE = 16'h1296;
		1954: SAMPLE = 16'h1264;
		1955: SAMPLE = 16'h1232;
		1956: SAMPLE = 16'h1201;
		1957: SAMPLE = 16'h11cf;
		1958: SAMPLE = 16'h119d;
		1959: SAMPLE = 16'h116b;
		1960: SAMPLE = 16'h1139;
		1961: SAMPLE = 16'h1108;
		1962: SAMPLE = 16'h10d6;
		1963: SAMPLE = 16'h10a4;
		1964: SAMPLE = 16'h1072;
		1965: SAMPLE = 16'h1040;
		1966: SAMPLE = 16'h100e;
		1967: SAMPLE = 16'hfdd;
		1968: SAMPLE = 16'hfab;
		1969: SAMPLE = 16'hf79;
		1970: SAMPLE = 16'hf47;
		1971: SAMPLE = 16'hf15;
		1972: SAMPLE = 16'hee3;
		1973: SAMPLE = 16'heb1;
		1974: SAMPLE = 16'he7f;
		1975: SAMPLE = 16'he4d;
		1976: SAMPLE = 16'he1b;
		1977: SAMPLE = 16'hde9;
		1978: SAMPLE = 16'hdb7;
		1979: SAMPLE = 16'hd85;
		1980: SAMPLE = 16'hd53;
		1981: SAMPLE = 16'hd21;
		1982: SAMPLE = 16'hcef;
		1983: SAMPLE = 16'hcbd;
		1984: SAMPLE = 16'hc8b;
		1985: SAMPLE = 16'hc59;
		1986: SAMPLE = 16'hc27;
		1987: SAMPLE = 16'hbf5;
		1988: SAMPLE = 16'hbc3;
		1989: SAMPLE = 16'hb91;
		1990: SAMPLE = 16'hb5f;
		1991: SAMPLE = 16'hb2d;
		1992: SAMPLE = 16'hafb;
		1993: SAMPLE = 16'hac9;
		1994: SAMPLE = 16'ha97;
		1995: SAMPLE = 16'ha65;
		1996: SAMPLE = 16'ha33;
		1997: SAMPLE = 16'ha00;
		1998: SAMPLE = 16'h9ce;
		1999: SAMPLE = 16'h99c;
		2000: SAMPLE = 16'h96a;
		2001: SAMPLE = 16'h938;
		2002: SAMPLE = 16'h906;
		2003: SAMPLE = 16'h8d4;
		2004: SAMPLE = 16'h8a2;
		2005: SAMPLE = 16'h86f;
		2006: SAMPLE = 16'h83d;
		2007: SAMPLE = 16'h80b;
		2008: SAMPLE = 16'h7d9;
		2009: SAMPLE = 16'h7a7;
		2010: SAMPLE = 16'h775;
		2011: SAMPLE = 16'h742;
		2012: SAMPLE = 16'h710;
		2013: SAMPLE = 16'h6de;
		2014: SAMPLE = 16'h6ac;
		2015: SAMPLE = 16'h67a;
		2016: SAMPLE = 16'h647;
		2017: SAMPLE = 16'h615;
		2018: SAMPLE = 16'h5e3;
		2019: SAMPLE = 16'h5b1;
		2020: SAMPLE = 16'h57f;
		2021: SAMPLE = 16'h54c;
		2022: SAMPLE = 16'h51a;
		2023: SAMPLE = 16'h4e8;
		2024: SAMPLE = 16'h4b6;
		2025: SAMPLE = 16'h483;
		2026: SAMPLE = 16'h451;
		2027: SAMPLE = 16'h41f;
		2028: SAMPLE = 16'h3ed;
		2029: SAMPLE = 16'h3ba;
		2030: SAMPLE = 16'h388;
		2031: SAMPLE = 16'h356;
		2032: SAMPLE = 16'h324;
		2033: SAMPLE = 16'h2f1;
		2034: SAMPLE = 16'h2bf;
		2035: SAMPLE = 16'h28d;
		2036: SAMPLE = 16'h25b;
		2037: SAMPLE = 16'h228;
		2038: SAMPLE = 16'h1f6;
		2039: SAMPLE = 16'h1c4;
		2040: SAMPLE = 16'h192;
		2041: SAMPLE = 16'h15f;
		2042: SAMPLE = 16'h12d;
		2043: SAMPLE = 16'hfb;
		2044: SAMPLE = 16'hc9;
		2045: SAMPLE = 16'h96;
		2046: SAMPLE = 16'h64;
		2047: SAMPLE = 16'h32;
		2048: SAMPLE = 16'h0;
		2049: SAMPLE = 16'hffcd;
		2050: SAMPLE = 16'hff9b;
		2051: SAMPLE = 16'hff69;
		2052: SAMPLE = 16'hff36;
		2053: SAMPLE = 16'hff04;
		2054: SAMPLE = 16'hfed2;
		2055: SAMPLE = 16'hfea0;
		2056: SAMPLE = 16'hfe6d;
		2057: SAMPLE = 16'hfe3b;
		2058: SAMPLE = 16'hfe09;
		2059: SAMPLE = 16'hfdd7;
		2060: SAMPLE = 16'hfda4;
		2061: SAMPLE = 16'hfd72;
		2062: SAMPLE = 16'hfd40;
		2063: SAMPLE = 16'hfd0e;
		2064: SAMPLE = 16'hfcdb;
		2065: SAMPLE = 16'hfca9;
		2066: SAMPLE = 16'hfc77;
		2067: SAMPLE = 16'hfc45;
		2068: SAMPLE = 16'hfc12;
		2069: SAMPLE = 16'hfbe0;
		2070: SAMPLE = 16'hfbae;
		2071: SAMPLE = 16'hfb7c;
		2072: SAMPLE = 16'hfb49;
		2073: SAMPLE = 16'hfb17;
		2074: SAMPLE = 16'hfae5;
		2075: SAMPLE = 16'hfab3;
		2076: SAMPLE = 16'hfa80;
		2077: SAMPLE = 16'hfa4e;
		2078: SAMPLE = 16'hfa1c;
		2079: SAMPLE = 16'hf9ea;
		2080: SAMPLE = 16'hf9b8;
		2081: SAMPLE = 16'hf985;
		2082: SAMPLE = 16'hf953;
		2083: SAMPLE = 16'hf921;
		2084: SAMPLE = 16'hf8ef;
		2085: SAMPLE = 16'hf8bd;
		2086: SAMPLE = 16'hf88a;
		2087: SAMPLE = 16'hf858;
		2088: SAMPLE = 16'hf826;
		2089: SAMPLE = 16'hf7f4;
		2090: SAMPLE = 16'hf7c2;
		2091: SAMPLE = 16'hf790;
		2092: SAMPLE = 16'hf75d;
		2093: SAMPLE = 16'hf72b;
		2094: SAMPLE = 16'hf6f9;
		2095: SAMPLE = 16'hf6c7;
		2096: SAMPLE = 16'hf695;
		2097: SAMPLE = 16'hf663;
		2098: SAMPLE = 16'hf631;
		2099: SAMPLE = 16'hf5ff;
		2100: SAMPLE = 16'hf5cc;
		2101: SAMPLE = 16'hf59a;
		2102: SAMPLE = 16'hf568;
		2103: SAMPLE = 16'hf536;
		2104: SAMPLE = 16'hf504;
		2105: SAMPLE = 16'hf4d2;
		2106: SAMPLE = 16'hf4a0;
		2107: SAMPLE = 16'hf46e;
		2108: SAMPLE = 16'hf43c;
		2109: SAMPLE = 16'hf40a;
		2110: SAMPLE = 16'hf3d8;
		2111: SAMPLE = 16'hf3a6;
		2112: SAMPLE = 16'hf374;
		2113: SAMPLE = 16'hf342;
		2114: SAMPLE = 16'hf310;
		2115: SAMPLE = 16'hf2de;
		2116: SAMPLE = 16'hf2ac;
		2117: SAMPLE = 16'hf27a;
		2118: SAMPLE = 16'hf248;
		2119: SAMPLE = 16'hf216;
		2120: SAMPLE = 16'hf1e4;
		2121: SAMPLE = 16'hf1b2;
		2122: SAMPLE = 16'hf180;
		2123: SAMPLE = 16'hf14e;
		2124: SAMPLE = 16'hf11c;
		2125: SAMPLE = 16'hf0ea;
		2126: SAMPLE = 16'hf0b8;
		2127: SAMPLE = 16'hf086;
		2128: SAMPLE = 16'hf054;
		2129: SAMPLE = 16'hf022;
		2130: SAMPLE = 16'heff1;
		2131: SAMPLE = 16'hefbf;
		2132: SAMPLE = 16'hef8d;
		2133: SAMPLE = 16'hef5b;
		2134: SAMPLE = 16'hef29;
		2135: SAMPLE = 16'heef7;
		2136: SAMPLE = 16'heec6;
		2137: SAMPLE = 16'hee94;
		2138: SAMPLE = 16'hee62;
		2139: SAMPLE = 16'hee30;
		2140: SAMPLE = 16'hedfe;
		2141: SAMPLE = 16'hedcd;
		2142: SAMPLE = 16'hed9b;
		2143: SAMPLE = 16'hed69;
		2144: SAMPLE = 16'hed37;
		2145: SAMPLE = 16'hed06;
		2146: SAMPLE = 16'hecd4;
		2147: SAMPLE = 16'heca2;
		2148: SAMPLE = 16'hec71;
		2149: SAMPLE = 16'hec3f;
		2150: SAMPLE = 16'hec0d;
		2151: SAMPLE = 16'hebdc;
		2152: SAMPLE = 16'hebaa;
		2153: SAMPLE = 16'heb78;
		2154: SAMPLE = 16'heb47;
		2155: SAMPLE = 16'heb15;
		2156: SAMPLE = 16'heae4;
		2157: SAMPLE = 16'heab2;
		2158: SAMPLE = 16'hea80;
		2159: SAMPLE = 16'hea4f;
		2160: SAMPLE = 16'hea1d;
		2161: SAMPLE = 16'he9ec;
		2162: SAMPLE = 16'he9ba;
		2163: SAMPLE = 16'he989;
		2164: SAMPLE = 16'he957;
		2165: SAMPLE = 16'he926;
		2166: SAMPLE = 16'he8f5;
		2167: SAMPLE = 16'he8c3;
		2168: SAMPLE = 16'he892;
		2169: SAMPLE = 16'he860;
		2170: SAMPLE = 16'he82f;
		2171: SAMPLE = 16'he7fd;
		2172: SAMPLE = 16'he7cc;
		2173: SAMPLE = 16'he79b;
		2174: SAMPLE = 16'he769;
		2175: SAMPLE = 16'he738;
		2176: SAMPLE = 16'he707;
		2177: SAMPLE = 16'he6d5;
		2178: SAMPLE = 16'he6a4;
		2179: SAMPLE = 16'he673;
		2180: SAMPLE = 16'he642;
		2181: SAMPLE = 16'he610;
		2182: SAMPLE = 16'he5df;
		2183: SAMPLE = 16'he5ae;
		2184: SAMPLE = 16'he57d;
		2185: SAMPLE = 16'he54c;
		2186: SAMPLE = 16'he51b;
		2187: SAMPLE = 16'he4e9;
		2188: SAMPLE = 16'he4b8;
		2189: SAMPLE = 16'he487;
		2190: SAMPLE = 16'he456;
		2191: SAMPLE = 16'he425;
		2192: SAMPLE = 16'he3f4;
		2193: SAMPLE = 16'he3c3;
		2194: SAMPLE = 16'he392;
		2195: SAMPLE = 16'he361;
		2196: SAMPLE = 16'he330;
		2197: SAMPLE = 16'he2ff;
		2198: SAMPLE = 16'he2ce;
		2199: SAMPLE = 16'he29d;
		2200: SAMPLE = 16'he26c;
		2201: SAMPLE = 16'he23b;
		2202: SAMPLE = 16'he20a;
		2203: SAMPLE = 16'he1da;
		2204: SAMPLE = 16'he1a9;
		2205: SAMPLE = 16'he178;
		2206: SAMPLE = 16'he147;
		2207: SAMPLE = 16'he116;
		2208: SAMPLE = 16'he0e6;
		2209: SAMPLE = 16'he0b5;
		2210: SAMPLE = 16'he084;
		2211: SAMPLE = 16'he053;
		2212: SAMPLE = 16'he023;
		2213: SAMPLE = 16'hdff2;
		2214: SAMPLE = 16'hdfc1;
		2215: SAMPLE = 16'hdf91;
		2216: SAMPLE = 16'hdf60;
		2217: SAMPLE = 16'hdf2f;
		2218: SAMPLE = 16'hdeff;
		2219: SAMPLE = 16'hdece;
		2220: SAMPLE = 16'hde9e;
		2221: SAMPLE = 16'hde6d;
		2222: SAMPLE = 16'hde3d;
		2223: SAMPLE = 16'hde0c;
		2224: SAMPLE = 16'hdddc;
		2225: SAMPLE = 16'hddab;
		2226: SAMPLE = 16'hdd7b;
		2227: SAMPLE = 16'hdd4b;
		2228: SAMPLE = 16'hdd1a;
		2229: SAMPLE = 16'hdcea;
		2230: SAMPLE = 16'hdcba;
		2231: SAMPLE = 16'hdc89;
		2232: SAMPLE = 16'hdc59;
		2233: SAMPLE = 16'hdc29;
		2234: SAMPLE = 16'hdbf8;
		2235: SAMPLE = 16'hdbc8;
		2236: SAMPLE = 16'hdb98;
		2237: SAMPLE = 16'hdb68;
		2238: SAMPLE = 16'hdb38;
		2239: SAMPLE = 16'hdb08;
		2240: SAMPLE = 16'hdad7;
		2241: SAMPLE = 16'hdaa7;
		2242: SAMPLE = 16'hda77;
		2243: SAMPLE = 16'hda47;
		2244: SAMPLE = 16'hda17;
		2245: SAMPLE = 16'hd9e7;
		2246: SAMPLE = 16'hd9b7;
		2247: SAMPLE = 16'hd987;
		2248: SAMPLE = 16'hd957;
		2249: SAMPLE = 16'hd927;
		2250: SAMPLE = 16'hd8f8;
		2251: SAMPLE = 16'hd8c8;
		2252: SAMPLE = 16'hd898;
		2253: SAMPLE = 16'hd868;
		2254: SAMPLE = 16'hd838;
		2255: SAMPLE = 16'hd809;
		2256: SAMPLE = 16'hd7d9;
		2257: SAMPLE = 16'hd7a9;
		2258: SAMPLE = 16'hd779;
		2259: SAMPLE = 16'hd74a;
		2260: SAMPLE = 16'hd71a;
		2261: SAMPLE = 16'hd6ea;
		2262: SAMPLE = 16'hd6bb;
		2263: SAMPLE = 16'hd68b;
		2264: SAMPLE = 16'hd65c;
		2265: SAMPLE = 16'hd62c;
		2266: SAMPLE = 16'hd5fd;
		2267: SAMPLE = 16'hd5cd;
		2268: SAMPLE = 16'hd59e;
		2269: SAMPLE = 16'hd56e;
		2270: SAMPLE = 16'hd53f;
		2271: SAMPLE = 16'hd510;
		2272: SAMPLE = 16'hd4e0;
		2273: SAMPLE = 16'hd4b1;
		2274: SAMPLE = 16'hd482;
		2275: SAMPLE = 16'hd452;
		2276: SAMPLE = 16'hd423;
		2277: SAMPLE = 16'hd3f4;
		2278: SAMPLE = 16'hd3c5;
		2279: SAMPLE = 16'hd396;
		2280: SAMPLE = 16'hd367;
		2281: SAMPLE = 16'hd337;
		2282: SAMPLE = 16'hd308;
		2283: SAMPLE = 16'hd2d9;
		2284: SAMPLE = 16'hd2aa;
		2285: SAMPLE = 16'hd27b;
		2286: SAMPLE = 16'hd24c;
		2287: SAMPLE = 16'hd21d;
		2288: SAMPLE = 16'hd1ee;
		2289: SAMPLE = 16'hd1c0;
		2290: SAMPLE = 16'hd191;
		2291: SAMPLE = 16'hd162;
		2292: SAMPLE = 16'hd133;
		2293: SAMPLE = 16'hd104;
		2294: SAMPLE = 16'hd0d6;
		2295: SAMPLE = 16'hd0a7;
		2296: SAMPLE = 16'hd078;
		2297: SAMPLE = 16'hd04a;
		2298: SAMPLE = 16'hd01b;
		2299: SAMPLE = 16'hcfec;
		2300: SAMPLE = 16'hcfbe;
		2301: SAMPLE = 16'hcf8f;
		2302: SAMPLE = 16'hcf61;
		2303: SAMPLE = 16'hcf32;
		2304: SAMPLE = 16'hcf04;
		2305: SAMPLE = 16'hced5;
		2306: SAMPLE = 16'hcea7;
		2307: SAMPLE = 16'hce79;
		2308: SAMPLE = 16'hce4a;
		2309: SAMPLE = 16'hce1c;
		2310: SAMPLE = 16'hcdee;
		2311: SAMPLE = 16'hcdbf;
		2312: SAMPLE = 16'hcd91;
		2313: SAMPLE = 16'hcd63;
		2314: SAMPLE = 16'hcd35;
		2315: SAMPLE = 16'hcd07;
		2316: SAMPLE = 16'hccd9;
		2317: SAMPLE = 16'hccab;
		2318: SAMPLE = 16'hcc7d;
		2319: SAMPLE = 16'hcc4f;
		2320: SAMPLE = 16'hcc21;
		2321: SAMPLE = 16'hcbf3;
		2322: SAMPLE = 16'hcbc5;
		2323: SAMPLE = 16'hcb97;
		2324: SAMPLE = 16'hcb69;
		2325: SAMPLE = 16'hcb3b;
		2326: SAMPLE = 16'hcb0d;
		2327: SAMPLE = 16'hcae0;
		2328: SAMPLE = 16'hcab2;
		2329: SAMPLE = 16'hca84;
		2330: SAMPLE = 16'hca57;
		2331: SAMPLE = 16'hca29;
		2332: SAMPLE = 16'hc9fb;
		2333: SAMPLE = 16'hc9ce;
		2334: SAMPLE = 16'hc9a0;
		2335: SAMPLE = 16'hc973;
		2336: SAMPLE = 16'hc945;
		2337: SAMPLE = 16'hc918;
		2338: SAMPLE = 16'hc8eb;
		2339: SAMPLE = 16'hc8bd;
		2340: SAMPLE = 16'hc890;
		2341: SAMPLE = 16'hc863;
		2342: SAMPLE = 16'hc835;
		2343: SAMPLE = 16'hc808;
		2344: SAMPLE = 16'hc7db;
		2345: SAMPLE = 16'hc7ae;
		2346: SAMPLE = 16'hc781;
		2347: SAMPLE = 16'hc754;
		2348: SAMPLE = 16'hc727;
		2349: SAMPLE = 16'hc6f9;
		2350: SAMPLE = 16'hc6cd;
		2351: SAMPLE = 16'hc6a0;
		2352: SAMPLE = 16'hc673;
		2353: SAMPLE = 16'hc646;
		2354: SAMPLE = 16'hc619;
		2355: SAMPLE = 16'hc5ec;
		2356: SAMPLE = 16'hc5bf;
		2357: SAMPLE = 16'hc593;
		2358: SAMPLE = 16'hc566;
		2359: SAMPLE = 16'hc539;
		2360: SAMPLE = 16'hc50d;
		2361: SAMPLE = 16'hc4e0;
		2362: SAMPLE = 16'hc4b3;
		2363: SAMPLE = 16'hc487;
		2364: SAMPLE = 16'hc45a;
		2365: SAMPLE = 16'hc42e;
		2366: SAMPLE = 16'hc402;
		2367: SAMPLE = 16'hc3d5;
		2368: SAMPLE = 16'hc3a9;
		2369: SAMPLE = 16'hc37c;
		2370: SAMPLE = 16'hc350;
		2371: SAMPLE = 16'hc324;
		2372: SAMPLE = 16'hc2f8;
		2373: SAMPLE = 16'hc2cc;
		2374: SAMPLE = 16'hc29f;
		2375: SAMPLE = 16'hc273;
		2376: SAMPLE = 16'hc247;
		2377: SAMPLE = 16'hc21b;
		2378: SAMPLE = 16'hc1ef;
		2379: SAMPLE = 16'hc1c3;
		2380: SAMPLE = 16'hc197;
		2381: SAMPLE = 16'hc16c;
		2382: SAMPLE = 16'hc140;
		2383: SAMPLE = 16'hc114;
		2384: SAMPLE = 16'hc0e8;
		2385: SAMPLE = 16'hc0bc;
		2386: SAMPLE = 16'hc091;
		2387: SAMPLE = 16'hc065;
		2388: SAMPLE = 16'hc03a;
		2389: SAMPLE = 16'hc00e;
		2390: SAMPLE = 16'hbfe2;
		2391: SAMPLE = 16'hbfb7;
		2392: SAMPLE = 16'hbf8c;
		2393: SAMPLE = 16'hbf60;
		2394: SAMPLE = 16'hbf35;
		2395: SAMPLE = 16'hbf09;
		2396: SAMPLE = 16'hbede;
		2397: SAMPLE = 16'hbeb3;
		2398: SAMPLE = 16'hbe88;
		2399: SAMPLE = 16'hbe5d;
		2400: SAMPLE = 16'hbe31;
		2401: SAMPLE = 16'hbe06;
		2402: SAMPLE = 16'hbddb;
		2403: SAMPLE = 16'hbdb0;
		2404: SAMPLE = 16'hbd85;
		2405: SAMPLE = 16'hbd5a;
		2406: SAMPLE = 16'hbd2f;
		2407: SAMPLE = 16'hbd05;
		2408: SAMPLE = 16'hbcda;
		2409: SAMPLE = 16'hbcaf;
		2410: SAMPLE = 16'hbc84;
		2411: SAMPLE = 16'hbc5a;
		2412: SAMPLE = 16'hbc2f;
		2413: SAMPLE = 16'hbc04;
		2414: SAMPLE = 16'hbbda;
		2415: SAMPLE = 16'hbbaf;
		2416: SAMPLE = 16'hbb85;
		2417: SAMPLE = 16'hbb5a;
		2418: SAMPLE = 16'hbb30;
		2419: SAMPLE = 16'hbb05;
		2420: SAMPLE = 16'hbadb;
		2421: SAMPLE = 16'hbab1;
		2422: SAMPLE = 16'hba87;
		2423: SAMPLE = 16'hba5c;
		2424: SAMPLE = 16'hba32;
		2425: SAMPLE = 16'hba08;
		2426: SAMPLE = 16'hb9de;
		2427: SAMPLE = 16'hb9b4;
		2428: SAMPLE = 16'hb98a;
		2429: SAMPLE = 16'hb960;
		2430: SAMPLE = 16'hb936;
		2431: SAMPLE = 16'hb90c;
		2432: SAMPLE = 16'hb8e3;
		2433: SAMPLE = 16'hb8b9;
		2434: SAMPLE = 16'hb88f;
		2435: SAMPLE = 16'hb865;
		2436: SAMPLE = 16'hb83c;
		2437: SAMPLE = 16'hb812;
		2438: SAMPLE = 16'hb7e9;
		2439: SAMPLE = 16'hb7bf;
		2440: SAMPLE = 16'hb796;
		2441: SAMPLE = 16'hb76c;
		2442: SAMPLE = 16'hb743;
		2443: SAMPLE = 16'hb719;
		2444: SAMPLE = 16'hb6f0;
		2445: SAMPLE = 16'hb6c7;
		2446: SAMPLE = 16'hb69e;
		2447: SAMPLE = 16'hb675;
		2448: SAMPLE = 16'hb64b;
		2449: SAMPLE = 16'hb622;
		2450: SAMPLE = 16'hb5f9;
		2451: SAMPLE = 16'hb5d0;
		2452: SAMPLE = 16'hb5a7;
		2453: SAMPLE = 16'hb57e;
		2454: SAMPLE = 16'hb556;
		2455: SAMPLE = 16'hb52d;
		2456: SAMPLE = 16'hb504;
		2457: SAMPLE = 16'hb4db;
		2458: SAMPLE = 16'hb4b3;
		2459: SAMPLE = 16'hb48a;
		2460: SAMPLE = 16'hb461;
		2461: SAMPLE = 16'hb439;
		2462: SAMPLE = 16'hb410;
		2463: SAMPLE = 16'hb3e8;
		2464: SAMPLE = 16'hb3c0;
		2465: SAMPLE = 16'hb397;
		2466: SAMPLE = 16'hb36f;
		2467: SAMPLE = 16'hb347;
		2468: SAMPLE = 16'hb31e;
		2469: SAMPLE = 16'hb2f6;
		2470: SAMPLE = 16'hb2ce;
		2471: SAMPLE = 16'hb2a6;
		2472: SAMPLE = 16'hb27e;
		2473: SAMPLE = 16'hb256;
		2474: SAMPLE = 16'hb22e;
		2475: SAMPLE = 16'hb206;
		2476: SAMPLE = 16'hb1de;
		2477: SAMPLE = 16'hb1b7;
		2478: SAMPLE = 16'hb18f;
		2479: SAMPLE = 16'hb167;
		2480: SAMPLE = 16'hb140;
		2481: SAMPLE = 16'hb118;
		2482: SAMPLE = 16'hb0f0;
		2483: SAMPLE = 16'hb0c9;
		2484: SAMPLE = 16'hb0a1;
		2485: SAMPLE = 16'hb07a;
		2486: SAMPLE = 16'hb053;
		2487: SAMPLE = 16'hb02b;
		2488: SAMPLE = 16'hb004;
		2489: SAMPLE = 16'hafdd;
		2490: SAMPLE = 16'hafb6;
		2491: SAMPLE = 16'haf8f;
		2492: SAMPLE = 16'haf68;
		2493: SAMPLE = 16'haf40;
		2494: SAMPLE = 16'haf1a;
		2495: SAMPLE = 16'haef3;
		2496: SAMPLE = 16'haecc;
		2497: SAMPLE = 16'haea5;
		2498: SAMPLE = 16'hae7e;
		2499: SAMPLE = 16'hae57;
		2500: SAMPLE = 16'hae31;
		2501: SAMPLE = 16'hae0a;
		2502: SAMPLE = 16'hade3;
		2503: SAMPLE = 16'hadbd;
		2504: SAMPLE = 16'had96;
		2505: SAMPLE = 16'had70;
		2506: SAMPLE = 16'had4a;
		2507: SAMPLE = 16'had23;
		2508: SAMPLE = 16'hacfd;
		2509: SAMPLE = 16'hacd7;
		2510: SAMPLE = 16'hacb1;
		2511: SAMPLE = 16'hac8a;
		2512: SAMPLE = 16'hac64;
		2513: SAMPLE = 16'hac3e;
		2514: SAMPLE = 16'hac18;
		2515: SAMPLE = 16'habf2;
		2516: SAMPLE = 16'habcc;
		2517: SAMPLE = 16'haba7;
		2518: SAMPLE = 16'hab81;
		2519: SAMPLE = 16'hab5b;
		2520: SAMPLE = 16'hab35;
		2521: SAMPLE = 16'hab10;
		2522: SAMPLE = 16'haaea;
		2523: SAMPLE = 16'haac5;
		2524: SAMPLE = 16'haa9f;
		2525: SAMPLE = 16'haa7a;
		2526: SAMPLE = 16'haa54;
		2527: SAMPLE = 16'haa2f;
		2528: SAMPLE = 16'haa0a;
		2529: SAMPLE = 16'ha9e5;
		2530: SAMPLE = 16'ha9bf;
		2531: SAMPLE = 16'ha99a;
		2532: SAMPLE = 16'ha975;
		2533: SAMPLE = 16'ha950;
		2534: SAMPLE = 16'ha92b;
		2535: SAMPLE = 16'ha906;
		2536: SAMPLE = 16'ha8e2;
		2537: SAMPLE = 16'ha8bd;
		2538: SAMPLE = 16'ha898;
		2539: SAMPLE = 16'ha873;
		2540: SAMPLE = 16'ha84f;
		2541: SAMPLE = 16'ha82a;
		2542: SAMPLE = 16'ha806;
		2543: SAMPLE = 16'ha7e1;
		2544: SAMPLE = 16'ha7bd;
		2545: SAMPLE = 16'ha798;
		2546: SAMPLE = 16'ha774;
		2547: SAMPLE = 16'ha750;
		2548: SAMPLE = 16'ha72b;
		2549: SAMPLE = 16'ha707;
		2550: SAMPLE = 16'ha6e3;
		2551: SAMPLE = 16'ha6bf;
		2552: SAMPLE = 16'ha69b;
		2553: SAMPLE = 16'ha677;
		2554: SAMPLE = 16'ha653;
		2555: SAMPLE = 16'ha62f;
		2556: SAMPLE = 16'ha60c;
		2557: SAMPLE = 16'ha5e8;
		2558: SAMPLE = 16'ha5c4;
		2559: SAMPLE = 16'ha5a1;
		2560: SAMPLE = 16'ha57d;
		2561: SAMPLE = 16'ha55a;
		2562: SAMPLE = 16'ha536;
		2563: SAMPLE = 16'ha513;
		2564: SAMPLE = 16'ha4ef;
		2565: SAMPLE = 16'ha4cc;
		2566: SAMPLE = 16'ha4a9;
		2567: SAMPLE = 16'ha486;
		2568: SAMPLE = 16'ha462;
		2569: SAMPLE = 16'ha43f;
		2570: SAMPLE = 16'ha41c;
		2571: SAMPLE = 16'ha3f9;
		2572: SAMPLE = 16'ha3d6;
		2573: SAMPLE = 16'ha3b4;
		2574: SAMPLE = 16'ha391;
		2575: SAMPLE = 16'ha36e;
		2576: SAMPLE = 16'ha34b;
		2577: SAMPLE = 16'ha329;
		2578: SAMPLE = 16'ha306;
		2579: SAMPLE = 16'ha2e4;
		2580: SAMPLE = 16'ha2c1;
		2581: SAMPLE = 16'ha29f;
		2582: SAMPLE = 16'ha27c;
		2583: SAMPLE = 16'ha25a;
		2584: SAMPLE = 16'ha238;
		2585: SAMPLE = 16'ha216;
		2586: SAMPLE = 16'ha1f4;
		2587: SAMPLE = 16'ha1d2;
		2588: SAMPLE = 16'ha1af;
		2589: SAMPLE = 16'ha18e;
		2590: SAMPLE = 16'ha16c;
		2591: SAMPLE = 16'ha14a;
		2592: SAMPLE = 16'ha128;
		2593: SAMPLE = 16'ha106;
		2594: SAMPLE = 16'ha0e5;
		2595: SAMPLE = 16'ha0c3;
		2596: SAMPLE = 16'ha0a1;
		2597: SAMPLE = 16'ha080;
		2598: SAMPLE = 16'ha05f;
		2599: SAMPLE = 16'ha03d;
		2600: SAMPLE = 16'ha01c;
		2601: SAMPLE = 16'h9ffb;
		2602: SAMPLE = 16'h9fd9;
		2603: SAMPLE = 16'h9fb8;
		2604: SAMPLE = 16'h9f97;
		2605: SAMPLE = 16'h9f76;
		2606: SAMPLE = 16'h9f55;
		2607: SAMPLE = 16'h9f34;
		2608: SAMPLE = 16'h9f13;
		2609: SAMPLE = 16'h9ef2;
		2610: SAMPLE = 16'h9ed2;
		2611: SAMPLE = 16'h9eb1;
		2612: SAMPLE = 16'h9e90;
		2613: SAMPLE = 16'h9e70;
		2614: SAMPLE = 16'h9e4f;
		2615: SAMPLE = 16'h9e2f;
		2616: SAMPLE = 16'h9e0e;
		2617: SAMPLE = 16'h9dee;
		2618: SAMPLE = 16'h9dce;
		2619: SAMPLE = 16'h9dae;
		2620: SAMPLE = 16'h9d8e;
		2621: SAMPLE = 16'h9d6d;
		2622: SAMPLE = 16'h9d4d;
		2623: SAMPLE = 16'h9d2d;
		2624: SAMPLE = 16'h9d0d;
		2625: SAMPLE = 16'h9cee;
		2626: SAMPLE = 16'h9cce;
		2627: SAMPLE = 16'h9cae;
		2628: SAMPLE = 16'h9c8e;
		2629: SAMPLE = 16'h9c6f;
		2630: SAMPLE = 16'h9c4f;
		2631: SAMPLE = 16'h9c30;
		2632: SAMPLE = 16'h9c10;
		2633: SAMPLE = 16'h9bf1;
		2634: SAMPLE = 16'h9bd2;
		2635: SAMPLE = 16'h9bb2;
		2636: SAMPLE = 16'h9b93;
		2637: SAMPLE = 16'h9b74;
		2638: SAMPLE = 16'h9b55;
		2639: SAMPLE = 16'h9b36;
		2640: SAMPLE = 16'h9b17;
		2641: SAMPLE = 16'h9af8;
		2642: SAMPLE = 16'h9ad9;
		2643: SAMPLE = 16'h9aba;
		2644: SAMPLE = 16'h9a9c;
		2645: SAMPLE = 16'h9a7d;
		2646: SAMPLE = 16'h9a5f;
		2647: SAMPLE = 16'h9a40;
		2648: SAMPLE = 16'h9a22;
		2649: SAMPLE = 16'h9a03;
		2650: SAMPLE = 16'h99e5;
		2651: SAMPLE = 16'h99c6;
		2652: SAMPLE = 16'h99a8;
		2653: SAMPLE = 16'h998a;
		2654: SAMPLE = 16'h996c;
		2655: SAMPLE = 16'h994e;
		2656: SAMPLE = 16'h9930;
		2657: SAMPLE = 16'h9912;
		2658: SAMPLE = 16'h98f4;
		2659: SAMPLE = 16'h98d6;
		2660: SAMPLE = 16'h98b9;
		2661: SAMPLE = 16'h989b;
		2662: SAMPLE = 16'h987d;
		2663: SAMPLE = 16'h9860;
		2664: SAMPLE = 16'h9842;
		2665: SAMPLE = 16'h9825;
		2666: SAMPLE = 16'h9808;
		2667: SAMPLE = 16'h97ea;
		2668: SAMPLE = 16'h97cd;
		2669: SAMPLE = 16'h97b0;
		2670: SAMPLE = 16'h9793;
		2671: SAMPLE = 16'h9776;
		2672: SAMPLE = 16'h9759;
		2673: SAMPLE = 16'h973c;
		2674: SAMPLE = 16'h971f;
		2675: SAMPLE = 16'h9702;
		2676: SAMPLE = 16'h96e6;
		2677: SAMPLE = 16'h96c9;
		2678: SAMPLE = 16'h96ac;
		2679: SAMPLE = 16'h9690;
		2680: SAMPLE = 16'h9673;
		2681: SAMPLE = 16'h9657;
		2682: SAMPLE = 16'h963b;
		2683: SAMPLE = 16'h961e;
		2684: SAMPLE = 16'h9602;
		2685: SAMPLE = 16'h95e6;
		2686: SAMPLE = 16'h95ca;
		2687: SAMPLE = 16'h95ae;
		2688: SAMPLE = 16'h9592;
		2689: SAMPLE = 16'h9576;
		2690: SAMPLE = 16'h955a;
		2691: SAMPLE = 16'h953e;
		2692: SAMPLE = 16'h9523;
		2693: SAMPLE = 16'h9507;
		2694: SAMPLE = 16'h94ec;
		2695: SAMPLE = 16'h94d0;
		2696: SAMPLE = 16'h94b5;
		2697: SAMPLE = 16'h9499;
		2698: SAMPLE = 16'h947e;
		2699: SAMPLE = 16'h9463;
		2700: SAMPLE = 16'h9447;
		2701: SAMPLE = 16'h942c;
		2702: SAMPLE = 16'h9411;
		2703: SAMPLE = 16'h93f6;
		2704: SAMPLE = 16'h93db;
		2705: SAMPLE = 16'h93c0;
		2706: SAMPLE = 16'h93a6;
		2707: SAMPLE = 16'h938b;
		2708: SAMPLE = 16'h9370;
		2709: SAMPLE = 16'h9356;
		2710: SAMPLE = 16'h933b;
		2711: SAMPLE = 16'h9321;
		2712: SAMPLE = 16'h9306;
		2713: SAMPLE = 16'h92ec;
		2714: SAMPLE = 16'h92d2;
		2715: SAMPLE = 16'h92b7;
		2716: SAMPLE = 16'h929d;
		2717: SAMPLE = 16'h9283;
		2718: SAMPLE = 16'h9269;
		2719: SAMPLE = 16'h924f;
		2720: SAMPLE = 16'h9235;
		2721: SAMPLE = 16'h921c;
		2722: SAMPLE = 16'h9202;
		2723: SAMPLE = 16'h91e8;
		2724: SAMPLE = 16'h91cf;
		2725: SAMPLE = 16'h91b5;
		2726: SAMPLE = 16'h919c;
		2727: SAMPLE = 16'h9182;
		2728: SAMPLE = 16'h9169;
		2729: SAMPLE = 16'h9150;
		2730: SAMPLE = 16'h9136;
		2731: SAMPLE = 16'h911d;
		2732: SAMPLE = 16'h9104;
		2733: SAMPLE = 16'h90eb;
		2734: SAMPLE = 16'h90d2;
		2735: SAMPLE = 16'h90b9;
		2736: SAMPLE = 16'h90a0;
		2737: SAMPLE = 16'h9088;
		2738: SAMPLE = 16'h906f;
		2739: SAMPLE = 16'h9056;
		2740: SAMPLE = 16'h903e;
		2741: SAMPLE = 16'h9025;
		2742: SAMPLE = 16'h900d;
		2743: SAMPLE = 16'h8ff5;
		2744: SAMPLE = 16'h8fdc;
		2745: SAMPLE = 16'h8fc4;
		2746: SAMPLE = 16'h8fac;
		2747: SAMPLE = 16'h8f94;
		2748: SAMPLE = 16'h8f7c;
		2749: SAMPLE = 16'h8f64;
		2750: SAMPLE = 16'h8f4c;
		2751: SAMPLE = 16'h8f34;
		2752: SAMPLE = 16'h8f1d;
		2753: SAMPLE = 16'h8f05;
		2754: SAMPLE = 16'h8eed;
		2755: SAMPLE = 16'h8ed6;
		2756: SAMPLE = 16'h8ebe;
		2757: SAMPLE = 16'h8ea7;
		2758: SAMPLE = 16'h8e90;
		2759: SAMPLE = 16'h8e79;
		2760: SAMPLE = 16'h8e61;
		2761: SAMPLE = 16'h8e4a;
		2762: SAMPLE = 16'h8e33;
		2763: SAMPLE = 16'h8e1c;
		2764: SAMPLE = 16'h8e05;
		2765: SAMPLE = 16'h8dee;
		2766: SAMPLE = 16'h8dd8;
		2767: SAMPLE = 16'h8dc1;
		2768: SAMPLE = 16'h8daa;
		2769: SAMPLE = 16'h8d94;
		2770: SAMPLE = 16'h8d7d;
		2771: SAMPLE = 16'h8d67;
		2772: SAMPLE = 16'h8d50;
		2773: SAMPLE = 16'h8d3a;
		2774: SAMPLE = 16'h8d24;
		2775: SAMPLE = 16'h8d0e;
		2776: SAMPLE = 16'h8cf8;
		2777: SAMPLE = 16'h8ce2;
		2778: SAMPLE = 16'h8ccc;
		2779: SAMPLE = 16'h8cb6;
		2780: SAMPLE = 16'h8ca0;
		2781: SAMPLE = 16'h8c8a;
		2782: SAMPLE = 16'h8c75;
		2783: SAMPLE = 16'h8c5f;
		2784: SAMPLE = 16'h8c4a;
		2785: SAMPLE = 16'h8c34;
		2786: SAMPLE = 16'h8c1f;
		2787: SAMPLE = 16'h8c09;
		2788: SAMPLE = 16'h8bf4;
		2789: SAMPLE = 16'h8bdf;
		2790: SAMPLE = 16'h8bca;
		2791: SAMPLE = 16'h8bb5;
		2792: SAMPLE = 16'h8ba0;
		2793: SAMPLE = 16'h8b8b;
		2794: SAMPLE = 16'h8b76;
		2795: SAMPLE = 16'h8b61;
		2796: SAMPLE = 16'h8b4d;
		2797: SAMPLE = 16'h8b38;
		2798: SAMPLE = 16'h8b24;
		2799: SAMPLE = 16'h8b0f;
		2800: SAMPLE = 16'h8afb;
		2801: SAMPLE = 16'h8ae6;
		2802: SAMPLE = 16'h8ad2;
		2803: SAMPLE = 16'h8abe;
		2804: SAMPLE = 16'h8aaa;
		2805: SAMPLE = 16'h8a96;
		2806: SAMPLE = 16'h8a82;
		2807: SAMPLE = 16'h8a6e;
		2808: SAMPLE = 16'h8a5a;
		2809: SAMPLE = 16'h8a46;
		2810: SAMPLE = 16'h8a33;
		2811: SAMPLE = 16'h8a1f;
		2812: SAMPLE = 16'h8a0b;
		2813: SAMPLE = 16'h89f8;
		2814: SAMPLE = 16'h89e4;
		2815: SAMPLE = 16'h89d1;
		2816: SAMPLE = 16'h89be;
		2817: SAMPLE = 16'h89ab;
		2818: SAMPLE = 16'h8997;
		2819: SAMPLE = 16'h8984;
		2820: SAMPLE = 16'h8971;
		2821: SAMPLE = 16'h895f;
		2822: SAMPLE = 16'h894c;
		2823: SAMPLE = 16'h8939;
		2824: SAMPLE = 16'h8926;
		2825: SAMPLE = 16'h8914;
		2826: SAMPLE = 16'h8901;
		2827: SAMPLE = 16'h88ef;
		2828: SAMPLE = 16'h88dc;
		2829: SAMPLE = 16'h88ca;
		2830: SAMPLE = 16'h88b8;
		2831: SAMPLE = 16'h88a5;
		2832: SAMPLE = 16'h8893;
		2833: SAMPLE = 16'h8881;
		2834: SAMPLE = 16'h886f;
		2835: SAMPLE = 16'h885d;
		2836: SAMPLE = 16'h884b;
		2837: SAMPLE = 16'h883a;
		2838: SAMPLE = 16'h8828;
		2839: SAMPLE = 16'h8816;
		2840: SAMPLE = 16'h8805;
		2841: SAMPLE = 16'h87f3;
		2842: SAMPLE = 16'h87e2;
		2843: SAMPLE = 16'h87d1;
		2844: SAMPLE = 16'h87bf;
		2845: SAMPLE = 16'h87ae;
		2846: SAMPLE = 16'h879d;
		2847: SAMPLE = 16'h878c;
		2848: SAMPLE = 16'h877b;
		2849: SAMPLE = 16'h876a;
		2850: SAMPLE = 16'h8759;
		2851: SAMPLE = 16'h8749;
		2852: SAMPLE = 16'h8738;
		2853: SAMPLE = 16'h8727;
		2854: SAMPLE = 16'h8717;
		2855: SAMPLE = 16'h8706;
		2856: SAMPLE = 16'h86f6;
		2857: SAMPLE = 16'h86e6;
		2858: SAMPLE = 16'h86d5;
		2859: SAMPLE = 16'h86c5;
		2860: SAMPLE = 16'h86b5;
		2861: SAMPLE = 16'h86a5;
		2862: SAMPLE = 16'h8695;
		2863: SAMPLE = 16'h8685;
		2864: SAMPLE = 16'h8675;
		2865: SAMPLE = 16'h8666;
		2866: SAMPLE = 16'h8656;
		2867: SAMPLE = 16'h8646;
		2868: SAMPLE = 16'h8637;
		2869: SAMPLE = 16'h8627;
		2870: SAMPLE = 16'h8618;
		2871: SAMPLE = 16'h8609;
		2872: SAMPLE = 16'h85fa;
		2873: SAMPLE = 16'h85ea;
		2874: SAMPLE = 16'h85db;
		2875: SAMPLE = 16'h85cc;
		2876: SAMPLE = 16'h85bd;
		2877: SAMPLE = 16'h85af;
		2878: SAMPLE = 16'h85a0;
		2879: SAMPLE = 16'h8591;
		2880: SAMPLE = 16'h8582;
		2881: SAMPLE = 16'h8574;
		2882: SAMPLE = 16'h8565;
		2883: SAMPLE = 16'h8557;
		2884: SAMPLE = 16'h8549;
		2885: SAMPLE = 16'h853a;
		2886: SAMPLE = 16'h852c;
		2887: SAMPLE = 16'h851e;
		2888: SAMPLE = 16'h8510;
		2889: SAMPLE = 16'h8502;
		2890: SAMPLE = 16'h84f4;
		2891: SAMPLE = 16'h84e6;
		2892: SAMPLE = 16'h84d9;
		2893: SAMPLE = 16'h84cb;
		2894: SAMPLE = 16'h84bd;
		2895: SAMPLE = 16'h84b0;
		2896: SAMPLE = 16'h84a2;
		2897: SAMPLE = 16'h8495;
		2898: SAMPLE = 16'h8488;
		2899: SAMPLE = 16'h847b;
		2900: SAMPLE = 16'h846d;
		2901: SAMPLE = 16'h8460;
		2902: SAMPLE = 16'h8453;
		2903: SAMPLE = 16'h8446;
		2904: SAMPLE = 16'h843a;
		2905: SAMPLE = 16'h842d;
		2906: SAMPLE = 16'h8420;
		2907: SAMPLE = 16'h8414;
		2908: SAMPLE = 16'h8407;
		2909: SAMPLE = 16'h83fa;
		2910: SAMPLE = 16'h83ee;
		2911: SAMPLE = 16'h83e2;
		2912: SAMPLE = 16'h83d6;
		2913: SAMPLE = 16'h83c9;
		2914: SAMPLE = 16'h83bd;
		2915: SAMPLE = 16'h83b1;
		2916: SAMPLE = 16'h83a5;
		2917: SAMPLE = 16'h8399;
		2918: SAMPLE = 16'h838e;
		2919: SAMPLE = 16'h8382;
		2920: SAMPLE = 16'h8376;
		2921: SAMPLE = 16'h836b;
		2922: SAMPLE = 16'h835f;
		2923: SAMPLE = 16'h8354;
		2924: SAMPLE = 16'h8348;
		2925: SAMPLE = 16'h833d;
		2926: SAMPLE = 16'h8332;
		2927: SAMPLE = 16'h8327;
		2928: SAMPLE = 16'h831c;
		2929: SAMPLE = 16'h8311;
		2930: SAMPLE = 16'h8306;
		2931: SAMPLE = 16'h82fb;
		2932: SAMPLE = 16'h82f0;
		2933: SAMPLE = 16'h82e6;
		2934: SAMPLE = 16'h82db;
		2935: SAMPLE = 16'h82d0;
		2936: SAMPLE = 16'h82c6;
		2937: SAMPLE = 16'h82bc;
		2938: SAMPLE = 16'h82b1;
		2939: SAMPLE = 16'h82a7;
		2940: SAMPLE = 16'h829d;
		2941: SAMPLE = 16'h8293;
		2942: SAMPLE = 16'h8289;
		2943: SAMPLE = 16'h827f;
		2944: SAMPLE = 16'h8275;
		2945: SAMPLE = 16'h826b;
		2946: SAMPLE = 16'h8262;
		2947: SAMPLE = 16'h8258;
		2948: SAMPLE = 16'h824f;
		2949: SAMPLE = 16'h8245;
		2950: SAMPLE = 16'h823c;
		2951: SAMPLE = 16'h8232;
		2952: SAMPLE = 16'h8229;
		2953: SAMPLE = 16'h8220;
		2954: SAMPLE = 16'h8217;
		2955: SAMPLE = 16'h820e;
		2956: SAMPLE = 16'h8205;
		2957: SAMPLE = 16'h81fc;
		2958: SAMPLE = 16'h81f3;
		2959: SAMPLE = 16'h81eb;
		2960: SAMPLE = 16'h81e2;
		2961: SAMPLE = 16'h81d9;
		2962: SAMPLE = 16'h81d1;
		2963: SAMPLE = 16'h81c8;
		2964: SAMPLE = 16'h81c0;
		2965: SAMPLE = 16'h81b8;
		2966: SAMPLE = 16'h81b0;
		2967: SAMPLE = 16'h81a8;
		2968: SAMPLE = 16'h81a0;
		2969: SAMPLE = 16'h8198;
		2970: SAMPLE = 16'h8190;
		2971: SAMPLE = 16'h8188;
		2972: SAMPLE = 16'h8180;
		2973: SAMPLE = 16'h8179;
		2974: SAMPLE = 16'h8171;
		2975: SAMPLE = 16'h816a;
		2976: SAMPLE = 16'h8162;
		2977: SAMPLE = 16'h815b;
		2978: SAMPLE = 16'h8154;
		2979: SAMPLE = 16'h814c;
		2980: SAMPLE = 16'h8145;
		2981: SAMPLE = 16'h813e;
		2982: SAMPLE = 16'h8137;
		2983: SAMPLE = 16'h8130;
		2984: SAMPLE = 16'h812a;
		2985: SAMPLE = 16'h8123;
		2986: SAMPLE = 16'h811c;
		2987: SAMPLE = 16'h8116;
		2988: SAMPLE = 16'h810f;
		2989: SAMPLE = 16'h8109;
		2990: SAMPLE = 16'h8102;
		2991: SAMPLE = 16'h80fc;
		2992: SAMPLE = 16'h80f6;
		2993: SAMPLE = 16'h80f0;
		2994: SAMPLE = 16'h80ea;
		2995: SAMPLE = 16'h80e4;
		2996: SAMPLE = 16'h80de;
		2997: SAMPLE = 16'h80d8;
		2998: SAMPLE = 16'h80d2;
		2999: SAMPLE = 16'h80cd;
		3000: SAMPLE = 16'h80c7;
		3001: SAMPLE = 16'h80c2;
		3002: SAMPLE = 16'h80bc;
		3003: SAMPLE = 16'h80b7;
		3004: SAMPLE = 16'h80b2;
		3005: SAMPLE = 16'h80ac;
		3006: SAMPLE = 16'h80a7;
		3007: SAMPLE = 16'h80a2;
		3008: SAMPLE = 16'h809d;
		3009: SAMPLE = 16'h8098;
		3010: SAMPLE = 16'h8094;
		3011: SAMPLE = 16'h808f;
		3012: SAMPLE = 16'h808a;
		3013: SAMPLE = 16'h8086;
		3014: SAMPLE = 16'h8081;
		3015: SAMPLE = 16'h807d;
		3016: SAMPLE = 16'h8078;
		3017: SAMPLE = 16'h8074;
		3018: SAMPLE = 16'h8070;
		3019: SAMPLE = 16'h806c;
		3020: SAMPLE = 16'h8068;
		3021: SAMPLE = 16'h8064;
		3022: SAMPLE = 16'h8060;
		3023: SAMPLE = 16'h805c;
		3024: SAMPLE = 16'h8058;
		3025: SAMPLE = 16'h8055;
		3026: SAMPLE = 16'h8051;
		3027: SAMPLE = 16'h804e;
		3028: SAMPLE = 16'h804a;
		3029: SAMPLE = 16'h8047;
		3030: SAMPLE = 16'h8043;
		3031: SAMPLE = 16'h8040;
		3032: SAMPLE = 16'h803d;
		3033: SAMPLE = 16'h803a;
		3034: SAMPLE = 16'h8037;
		3035: SAMPLE = 16'h8034;
		3036: SAMPLE = 16'h8031;
		3037: SAMPLE = 16'h802f;
		3038: SAMPLE = 16'h802c;
		3039: SAMPLE = 16'h8029;
		3040: SAMPLE = 16'h8027;
		3041: SAMPLE = 16'h8025;
		3042: SAMPLE = 16'h8022;
		3043: SAMPLE = 16'h8020;
		3044: SAMPLE = 16'h801e;
		3045: SAMPLE = 16'h801c;
		3046: SAMPLE = 16'h801a;
		3047: SAMPLE = 16'h8018;
		3048: SAMPLE = 16'h8016;
		3049: SAMPLE = 16'h8014;
		3050: SAMPLE = 16'h8012;
		3051: SAMPLE = 16'h8011;
		3052: SAMPLE = 16'h800f;
		3053: SAMPLE = 16'h800d;
		3054: SAMPLE = 16'h800c;
		3055: SAMPLE = 16'h800b;
		3056: SAMPLE = 16'h8009;
		3057: SAMPLE = 16'h8008;
		3058: SAMPLE = 16'h8007;
		3059: SAMPLE = 16'h8006;
		3060: SAMPLE = 16'h8005;
		3061: SAMPLE = 16'h8004;
		3062: SAMPLE = 16'h8003;
		3063: SAMPLE = 16'h8003;
		3064: SAMPLE = 16'h8002;
		3065: SAMPLE = 16'h8001;
		3066: SAMPLE = 16'h8001;
		3067: SAMPLE = 16'h8000;
		3068: SAMPLE = 16'h8000;
		3069: SAMPLE = 16'h8000;
		3070: SAMPLE = 16'h8000;
		3071: SAMPLE = 16'h8000;
		3072: SAMPLE = 16'h8000;
		3073: SAMPLE = 16'h8000;
		3074: SAMPLE = 16'h8000;
		3075: SAMPLE = 16'h8000;
		3076: SAMPLE = 16'h8000;
		3077: SAMPLE = 16'h8000;
		3078: SAMPLE = 16'h8001;
		3079: SAMPLE = 16'h8001;
		3080: SAMPLE = 16'h8002;
		3081: SAMPLE = 16'h8003;
		3082: SAMPLE = 16'h8003;
		3083: SAMPLE = 16'h8004;
		3084: SAMPLE = 16'h8005;
		3085: SAMPLE = 16'h8006;
		3086: SAMPLE = 16'h8007;
		3087: SAMPLE = 16'h8008;
		3088: SAMPLE = 16'h8009;
		3089: SAMPLE = 16'h800b;
		3090: SAMPLE = 16'h800c;
		3091: SAMPLE = 16'h800d;
		3092: SAMPLE = 16'h800f;
		3093: SAMPLE = 16'h8011;
		3094: SAMPLE = 16'h8012;
		3095: SAMPLE = 16'h8014;
		3096: SAMPLE = 16'h8016;
		3097: SAMPLE = 16'h8018;
		3098: SAMPLE = 16'h801a;
		3099: SAMPLE = 16'h801c;
		3100: SAMPLE = 16'h801e;
		3101: SAMPLE = 16'h8020;
		3102: SAMPLE = 16'h8022;
		3103: SAMPLE = 16'h8025;
		3104: SAMPLE = 16'h8027;
		3105: SAMPLE = 16'h8029;
		3106: SAMPLE = 16'h802c;
		3107: SAMPLE = 16'h802f;
		3108: SAMPLE = 16'h8031;
		3109: SAMPLE = 16'h8034;
		3110: SAMPLE = 16'h8037;
		3111: SAMPLE = 16'h803a;
		3112: SAMPLE = 16'h803d;
		3113: SAMPLE = 16'h8040;
		3114: SAMPLE = 16'h8043;
		3115: SAMPLE = 16'h8047;
		3116: SAMPLE = 16'h804a;
		3117: SAMPLE = 16'h804e;
		3118: SAMPLE = 16'h8051;
		3119: SAMPLE = 16'h8055;
		3120: SAMPLE = 16'h8058;
		3121: SAMPLE = 16'h805c;
		3122: SAMPLE = 16'h8060;
		3123: SAMPLE = 16'h8064;
		3124: SAMPLE = 16'h8068;
		3125: SAMPLE = 16'h806c;
		3126: SAMPLE = 16'h8070;
		3127: SAMPLE = 16'h8074;
		3128: SAMPLE = 16'h8078;
		3129: SAMPLE = 16'h807d;
		3130: SAMPLE = 16'h8081;
		3131: SAMPLE = 16'h8086;
		3132: SAMPLE = 16'h808a;
		3133: SAMPLE = 16'h808f;
		3134: SAMPLE = 16'h8094;
		3135: SAMPLE = 16'h8098;
		3136: SAMPLE = 16'h809d;
		3137: SAMPLE = 16'h80a2;
		3138: SAMPLE = 16'h80a7;
		3139: SAMPLE = 16'h80ac;
		3140: SAMPLE = 16'h80b2;
		3141: SAMPLE = 16'h80b7;
		3142: SAMPLE = 16'h80bc;
		3143: SAMPLE = 16'h80c2;
		3144: SAMPLE = 16'h80c7;
		3145: SAMPLE = 16'h80cd;
		3146: SAMPLE = 16'h80d2;
		3147: SAMPLE = 16'h80d8;
		3148: SAMPLE = 16'h80de;
		3149: SAMPLE = 16'h80e4;
		3150: SAMPLE = 16'h80ea;
		3151: SAMPLE = 16'h80f0;
		3152: SAMPLE = 16'h80f6;
		3153: SAMPLE = 16'h80fc;
		3154: SAMPLE = 16'h8102;
		3155: SAMPLE = 16'h8109;
		3156: SAMPLE = 16'h810f;
		3157: SAMPLE = 16'h8116;
		3158: SAMPLE = 16'h811c;
		3159: SAMPLE = 16'h8123;
		3160: SAMPLE = 16'h812a;
		3161: SAMPLE = 16'h8130;
		3162: SAMPLE = 16'h8137;
		3163: SAMPLE = 16'h813e;
		3164: SAMPLE = 16'h8145;
		3165: SAMPLE = 16'h814c;
		3166: SAMPLE = 16'h8154;
		3167: SAMPLE = 16'h815b;
		3168: SAMPLE = 16'h8162;
		3169: SAMPLE = 16'h816a;
		3170: SAMPLE = 16'h8171;
		3171: SAMPLE = 16'h8179;
		3172: SAMPLE = 16'h8180;
		3173: SAMPLE = 16'h8188;
		3174: SAMPLE = 16'h8190;
		3175: SAMPLE = 16'h8198;
		3176: SAMPLE = 16'h81a0;
		3177: SAMPLE = 16'h81a8;
		3178: SAMPLE = 16'h81b0;
		3179: SAMPLE = 16'h81b8;
		3180: SAMPLE = 16'h81c0;
		3181: SAMPLE = 16'h81c8;
		3182: SAMPLE = 16'h81d1;
		3183: SAMPLE = 16'h81d9;
		3184: SAMPLE = 16'h81e2;
		3185: SAMPLE = 16'h81eb;
		3186: SAMPLE = 16'h81f3;
		3187: SAMPLE = 16'h81fc;
		3188: SAMPLE = 16'h8205;
		3189: SAMPLE = 16'h820e;
		3190: SAMPLE = 16'h8217;
		3191: SAMPLE = 16'h8220;
		3192: SAMPLE = 16'h8229;
		3193: SAMPLE = 16'h8232;
		3194: SAMPLE = 16'h823c;
		3195: SAMPLE = 16'h8245;
		3196: SAMPLE = 16'h824f;
		3197: SAMPLE = 16'h8258;
		3198: SAMPLE = 16'h8262;
		3199: SAMPLE = 16'h826b;
		3200: SAMPLE = 16'h8275;
		3201: SAMPLE = 16'h827f;
		3202: SAMPLE = 16'h8289;
		3203: SAMPLE = 16'h8293;
		3204: SAMPLE = 16'h829d;
		3205: SAMPLE = 16'h82a7;
		3206: SAMPLE = 16'h82b1;
		3207: SAMPLE = 16'h82bc;
		3208: SAMPLE = 16'h82c6;
		3209: SAMPLE = 16'h82d0;
		3210: SAMPLE = 16'h82db;
		3211: SAMPLE = 16'h82e6;
		3212: SAMPLE = 16'h82f0;
		3213: SAMPLE = 16'h82fb;
		3214: SAMPLE = 16'h8306;
		3215: SAMPLE = 16'h8311;
		3216: SAMPLE = 16'h831c;
		3217: SAMPLE = 16'h8327;
		3218: SAMPLE = 16'h8332;
		3219: SAMPLE = 16'h833d;
		3220: SAMPLE = 16'h8348;
		3221: SAMPLE = 16'h8354;
		3222: SAMPLE = 16'h835f;
		3223: SAMPLE = 16'h836b;
		3224: SAMPLE = 16'h8376;
		3225: SAMPLE = 16'h8382;
		3226: SAMPLE = 16'h838e;
		3227: SAMPLE = 16'h8399;
		3228: SAMPLE = 16'h83a5;
		3229: SAMPLE = 16'h83b1;
		3230: SAMPLE = 16'h83bd;
		3231: SAMPLE = 16'h83c9;
		3232: SAMPLE = 16'h83d6;
		3233: SAMPLE = 16'h83e2;
		3234: SAMPLE = 16'h83ee;
		3235: SAMPLE = 16'h83fa;
		3236: SAMPLE = 16'h8407;
		3237: SAMPLE = 16'h8414;
		3238: SAMPLE = 16'h8420;
		3239: SAMPLE = 16'h842d;
		3240: SAMPLE = 16'h843a;
		3241: SAMPLE = 16'h8446;
		3242: SAMPLE = 16'h8453;
		3243: SAMPLE = 16'h8460;
		3244: SAMPLE = 16'h846d;
		3245: SAMPLE = 16'h847b;
		3246: SAMPLE = 16'h8488;
		3247: SAMPLE = 16'h8495;
		3248: SAMPLE = 16'h84a2;
		3249: SAMPLE = 16'h84b0;
		3250: SAMPLE = 16'h84bd;
		3251: SAMPLE = 16'h84cb;
		3252: SAMPLE = 16'h84d9;
		3253: SAMPLE = 16'h84e6;
		3254: SAMPLE = 16'h84f4;
		3255: SAMPLE = 16'h8502;
		3256: SAMPLE = 16'h8510;
		3257: SAMPLE = 16'h851e;
		3258: SAMPLE = 16'h852c;
		3259: SAMPLE = 16'h853a;
		3260: SAMPLE = 16'h8549;
		3261: SAMPLE = 16'h8557;
		3262: SAMPLE = 16'h8565;
		3263: SAMPLE = 16'h8574;
		3264: SAMPLE = 16'h8582;
		3265: SAMPLE = 16'h8591;
		3266: SAMPLE = 16'h85a0;
		3267: SAMPLE = 16'h85af;
		3268: SAMPLE = 16'h85bd;
		3269: SAMPLE = 16'h85cc;
		3270: SAMPLE = 16'h85db;
		3271: SAMPLE = 16'h85ea;
		3272: SAMPLE = 16'h85fa;
		3273: SAMPLE = 16'h8609;
		3274: SAMPLE = 16'h8618;
		3275: SAMPLE = 16'h8627;
		3276: SAMPLE = 16'h8637;
		3277: SAMPLE = 16'h8646;
		3278: SAMPLE = 16'h8656;
		3279: SAMPLE = 16'h8666;
		3280: SAMPLE = 16'h8675;
		3281: SAMPLE = 16'h8685;
		3282: SAMPLE = 16'h8695;
		3283: SAMPLE = 16'h86a5;
		3284: SAMPLE = 16'h86b5;
		3285: SAMPLE = 16'h86c5;
		3286: SAMPLE = 16'h86d5;
		3287: SAMPLE = 16'h86e6;
		3288: SAMPLE = 16'h86f6;
		3289: SAMPLE = 16'h8706;
		3290: SAMPLE = 16'h8717;
		3291: SAMPLE = 16'h8727;
		3292: SAMPLE = 16'h8738;
		3293: SAMPLE = 16'h8749;
		3294: SAMPLE = 16'h8759;
		3295: SAMPLE = 16'h876a;
		3296: SAMPLE = 16'h877b;
		3297: SAMPLE = 16'h878c;
		3298: SAMPLE = 16'h879d;
		3299: SAMPLE = 16'h87ae;
		3300: SAMPLE = 16'h87bf;
		3301: SAMPLE = 16'h87d1;
		3302: SAMPLE = 16'h87e2;
		3303: SAMPLE = 16'h87f3;
		3304: SAMPLE = 16'h8805;
		3305: SAMPLE = 16'h8816;
		3306: SAMPLE = 16'h8828;
		3307: SAMPLE = 16'h883a;
		3308: SAMPLE = 16'h884b;
		3309: SAMPLE = 16'h885d;
		3310: SAMPLE = 16'h886f;
		3311: SAMPLE = 16'h8881;
		3312: SAMPLE = 16'h8893;
		3313: SAMPLE = 16'h88a5;
		3314: SAMPLE = 16'h88b8;
		3315: SAMPLE = 16'h88ca;
		3316: SAMPLE = 16'h88dc;
		3317: SAMPLE = 16'h88ef;
		3318: SAMPLE = 16'h8901;
		3319: SAMPLE = 16'h8914;
		3320: SAMPLE = 16'h8926;
		3321: SAMPLE = 16'h8939;
		3322: SAMPLE = 16'h894c;
		3323: SAMPLE = 16'h895f;
		3324: SAMPLE = 16'h8971;
		3325: SAMPLE = 16'h8984;
		3326: SAMPLE = 16'h8997;
		3327: SAMPLE = 16'h89ab;
		3328: SAMPLE = 16'h89be;
		3329: SAMPLE = 16'h89d1;
		3330: SAMPLE = 16'h89e4;
		3331: SAMPLE = 16'h89f8;
		3332: SAMPLE = 16'h8a0b;
		3333: SAMPLE = 16'h8a1f;
		3334: SAMPLE = 16'h8a33;
		3335: SAMPLE = 16'h8a46;
		3336: SAMPLE = 16'h8a5a;
		3337: SAMPLE = 16'h8a6e;
		3338: SAMPLE = 16'h8a82;
		3339: SAMPLE = 16'h8a96;
		3340: SAMPLE = 16'h8aaa;
		3341: SAMPLE = 16'h8abe;
		3342: SAMPLE = 16'h8ad2;
		3343: SAMPLE = 16'h8ae6;
		3344: SAMPLE = 16'h8afb;
		3345: SAMPLE = 16'h8b0f;
		3346: SAMPLE = 16'h8b24;
		3347: SAMPLE = 16'h8b38;
		3348: SAMPLE = 16'h8b4d;
		3349: SAMPLE = 16'h8b61;
		3350: SAMPLE = 16'h8b76;
		3351: SAMPLE = 16'h8b8b;
		3352: SAMPLE = 16'h8ba0;
		3353: SAMPLE = 16'h8bb5;
		3354: SAMPLE = 16'h8bca;
		3355: SAMPLE = 16'h8bdf;
		3356: SAMPLE = 16'h8bf4;
		3357: SAMPLE = 16'h8c09;
		3358: SAMPLE = 16'h8c1f;
		3359: SAMPLE = 16'h8c34;
		3360: SAMPLE = 16'h8c4a;
		3361: SAMPLE = 16'h8c5f;
		3362: SAMPLE = 16'h8c75;
		3363: SAMPLE = 16'h8c8a;
		3364: SAMPLE = 16'h8ca0;
		3365: SAMPLE = 16'h8cb6;
		3366: SAMPLE = 16'h8ccc;
		3367: SAMPLE = 16'h8ce2;
		3368: SAMPLE = 16'h8cf8;
		3369: SAMPLE = 16'h8d0e;
		3370: SAMPLE = 16'h8d24;
		3371: SAMPLE = 16'h8d3a;
		3372: SAMPLE = 16'h8d50;
		3373: SAMPLE = 16'h8d67;
		3374: SAMPLE = 16'h8d7d;
		3375: SAMPLE = 16'h8d94;
		3376: SAMPLE = 16'h8daa;
		3377: SAMPLE = 16'h8dc1;
		3378: SAMPLE = 16'h8dd8;
		3379: SAMPLE = 16'h8dee;
		3380: SAMPLE = 16'h8e05;
		3381: SAMPLE = 16'h8e1c;
		3382: SAMPLE = 16'h8e33;
		3383: SAMPLE = 16'h8e4a;
		3384: SAMPLE = 16'h8e61;
		3385: SAMPLE = 16'h8e79;
		3386: SAMPLE = 16'h8e90;
		3387: SAMPLE = 16'h8ea7;
		3388: SAMPLE = 16'h8ebe;
		3389: SAMPLE = 16'h8ed6;
		3390: SAMPLE = 16'h8eed;
		3391: SAMPLE = 16'h8f05;
		3392: SAMPLE = 16'h8f1d;
		3393: SAMPLE = 16'h8f34;
		3394: SAMPLE = 16'h8f4c;
		3395: SAMPLE = 16'h8f64;
		3396: SAMPLE = 16'h8f7c;
		3397: SAMPLE = 16'h8f94;
		3398: SAMPLE = 16'h8fac;
		3399: SAMPLE = 16'h8fc4;
		3400: SAMPLE = 16'h8fdc;
		3401: SAMPLE = 16'h8ff5;
		3402: SAMPLE = 16'h900d;
		3403: SAMPLE = 16'h9025;
		3404: SAMPLE = 16'h903e;
		3405: SAMPLE = 16'h9056;
		3406: SAMPLE = 16'h906f;
		3407: SAMPLE = 16'h9088;
		3408: SAMPLE = 16'h90a0;
		3409: SAMPLE = 16'h90b9;
		3410: SAMPLE = 16'h90d2;
		3411: SAMPLE = 16'h90eb;
		3412: SAMPLE = 16'h9104;
		3413: SAMPLE = 16'h911d;
		3414: SAMPLE = 16'h9136;
		3415: SAMPLE = 16'h9150;
		3416: SAMPLE = 16'h9169;
		3417: SAMPLE = 16'h9182;
		3418: SAMPLE = 16'h919c;
		3419: SAMPLE = 16'h91b5;
		3420: SAMPLE = 16'h91cf;
		3421: SAMPLE = 16'h91e8;
		3422: SAMPLE = 16'h9202;
		3423: SAMPLE = 16'h921c;
		3424: SAMPLE = 16'h9235;
		3425: SAMPLE = 16'h924f;
		3426: SAMPLE = 16'h9269;
		3427: SAMPLE = 16'h9283;
		3428: SAMPLE = 16'h929d;
		3429: SAMPLE = 16'h92b7;
		3430: SAMPLE = 16'h92d2;
		3431: SAMPLE = 16'h92ec;
		3432: SAMPLE = 16'h9306;
		3433: SAMPLE = 16'h9321;
		3434: SAMPLE = 16'h933b;
		3435: SAMPLE = 16'h9356;
		3436: SAMPLE = 16'h9370;
		3437: SAMPLE = 16'h938b;
		3438: SAMPLE = 16'h93a6;
		3439: SAMPLE = 16'h93c0;
		3440: SAMPLE = 16'h93db;
		3441: SAMPLE = 16'h93f6;
		3442: SAMPLE = 16'h9411;
		3443: SAMPLE = 16'h942c;
		3444: SAMPLE = 16'h9447;
		3445: SAMPLE = 16'h9463;
		3446: SAMPLE = 16'h947e;
		3447: SAMPLE = 16'h9499;
		3448: SAMPLE = 16'h94b5;
		3449: SAMPLE = 16'h94d0;
		3450: SAMPLE = 16'h94ec;
		3451: SAMPLE = 16'h9507;
		3452: SAMPLE = 16'h9523;
		3453: SAMPLE = 16'h953e;
		3454: SAMPLE = 16'h955a;
		3455: SAMPLE = 16'h9576;
		3456: SAMPLE = 16'h9592;
		3457: SAMPLE = 16'h95ae;
		3458: SAMPLE = 16'h95ca;
		3459: SAMPLE = 16'h95e6;
		3460: SAMPLE = 16'h9602;
		3461: SAMPLE = 16'h961e;
		3462: SAMPLE = 16'h963b;
		3463: SAMPLE = 16'h9657;
		3464: SAMPLE = 16'h9673;
		3465: SAMPLE = 16'h9690;
		3466: SAMPLE = 16'h96ac;
		3467: SAMPLE = 16'h96c9;
		3468: SAMPLE = 16'h96e6;
		3469: SAMPLE = 16'h9702;
		3470: SAMPLE = 16'h971f;
		3471: SAMPLE = 16'h973c;
		3472: SAMPLE = 16'h9759;
		3473: SAMPLE = 16'h9776;
		3474: SAMPLE = 16'h9793;
		3475: SAMPLE = 16'h97b0;
		3476: SAMPLE = 16'h97cd;
		3477: SAMPLE = 16'h97ea;
		3478: SAMPLE = 16'h9808;
		3479: SAMPLE = 16'h9825;
		3480: SAMPLE = 16'h9842;
		3481: SAMPLE = 16'h9860;
		3482: SAMPLE = 16'h987d;
		3483: SAMPLE = 16'h989b;
		3484: SAMPLE = 16'h98b9;
		3485: SAMPLE = 16'h98d6;
		3486: SAMPLE = 16'h98f4;
		3487: SAMPLE = 16'h9912;
		3488: SAMPLE = 16'h9930;
		3489: SAMPLE = 16'h994e;
		3490: SAMPLE = 16'h996c;
		3491: SAMPLE = 16'h998a;
		3492: SAMPLE = 16'h99a8;
		3493: SAMPLE = 16'h99c6;
		3494: SAMPLE = 16'h99e5;
		3495: SAMPLE = 16'h9a03;
		3496: SAMPLE = 16'h9a22;
		3497: SAMPLE = 16'h9a40;
		3498: SAMPLE = 16'h9a5f;
		3499: SAMPLE = 16'h9a7d;
		3500: SAMPLE = 16'h9a9c;
		3501: SAMPLE = 16'h9aba;
		3502: SAMPLE = 16'h9ad9;
		3503: SAMPLE = 16'h9af8;
		3504: SAMPLE = 16'h9b17;
		3505: SAMPLE = 16'h9b36;
		3506: SAMPLE = 16'h9b55;
		3507: SAMPLE = 16'h9b74;
		3508: SAMPLE = 16'h9b93;
		3509: SAMPLE = 16'h9bb2;
		3510: SAMPLE = 16'h9bd2;
		3511: SAMPLE = 16'h9bf1;
		3512: SAMPLE = 16'h9c10;
		3513: SAMPLE = 16'h9c30;
		3514: SAMPLE = 16'h9c4f;
		3515: SAMPLE = 16'h9c6f;
		3516: SAMPLE = 16'h9c8e;
		3517: SAMPLE = 16'h9cae;
		3518: SAMPLE = 16'h9cce;
		3519: SAMPLE = 16'h9cee;
		3520: SAMPLE = 16'h9d0d;
		3521: SAMPLE = 16'h9d2d;
		3522: SAMPLE = 16'h9d4d;
		3523: SAMPLE = 16'h9d6d;
		3524: SAMPLE = 16'h9d8e;
		3525: SAMPLE = 16'h9dae;
		3526: SAMPLE = 16'h9dce;
		3527: SAMPLE = 16'h9dee;
		3528: SAMPLE = 16'h9e0e;
		3529: SAMPLE = 16'h9e2f;
		3530: SAMPLE = 16'h9e4f;
		3531: SAMPLE = 16'h9e70;
		3532: SAMPLE = 16'h9e90;
		3533: SAMPLE = 16'h9eb1;
		3534: SAMPLE = 16'h9ed2;
		3535: SAMPLE = 16'h9ef2;
		3536: SAMPLE = 16'h9f13;
		3537: SAMPLE = 16'h9f34;
		3538: SAMPLE = 16'h9f55;
		3539: SAMPLE = 16'h9f76;
		3540: SAMPLE = 16'h9f97;
		3541: SAMPLE = 16'h9fb8;
		3542: SAMPLE = 16'h9fd9;
		3543: SAMPLE = 16'h9ffb;
		3544: SAMPLE = 16'ha01c;
		3545: SAMPLE = 16'ha03d;
		3546: SAMPLE = 16'ha05f;
		3547: SAMPLE = 16'ha080;
		3548: SAMPLE = 16'ha0a1;
		3549: SAMPLE = 16'ha0c3;
		3550: SAMPLE = 16'ha0e5;
		3551: SAMPLE = 16'ha106;
		3552: SAMPLE = 16'ha128;
		3553: SAMPLE = 16'ha14a;
		3554: SAMPLE = 16'ha16c;
		3555: SAMPLE = 16'ha18e;
		3556: SAMPLE = 16'ha1af;
		3557: SAMPLE = 16'ha1d2;
		3558: SAMPLE = 16'ha1f4;
		3559: SAMPLE = 16'ha216;
		3560: SAMPLE = 16'ha238;
		3561: SAMPLE = 16'ha25a;
		3562: SAMPLE = 16'ha27c;
		3563: SAMPLE = 16'ha29f;
		3564: SAMPLE = 16'ha2c1;
		3565: SAMPLE = 16'ha2e4;
		3566: SAMPLE = 16'ha306;
		3567: SAMPLE = 16'ha329;
		3568: SAMPLE = 16'ha34b;
		3569: SAMPLE = 16'ha36e;
		3570: SAMPLE = 16'ha391;
		3571: SAMPLE = 16'ha3b4;
		3572: SAMPLE = 16'ha3d6;
		3573: SAMPLE = 16'ha3f9;
		3574: SAMPLE = 16'ha41c;
		3575: SAMPLE = 16'ha43f;
		3576: SAMPLE = 16'ha462;
		3577: SAMPLE = 16'ha486;
		3578: SAMPLE = 16'ha4a9;
		3579: SAMPLE = 16'ha4cc;
		3580: SAMPLE = 16'ha4ef;
		3581: SAMPLE = 16'ha513;
		3582: SAMPLE = 16'ha536;
		3583: SAMPLE = 16'ha55a;
		3584: SAMPLE = 16'ha57d;
		3585: SAMPLE = 16'ha5a1;
		3586: SAMPLE = 16'ha5c4;
		3587: SAMPLE = 16'ha5e8;
		3588: SAMPLE = 16'ha60c;
		3589: SAMPLE = 16'ha62f;
		3590: SAMPLE = 16'ha653;
		3591: SAMPLE = 16'ha677;
		3592: SAMPLE = 16'ha69b;
		3593: SAMPLE = 16'ha6bf;
		3594: SAMPLE = 16'ha6e3;
		3595: SAMPLE = 16'ha707;
		3596: SAMPLE = 16'ha72b;
		3597: SAMPLE = 16'ha750;
		3598: SAMPLE = 16'ha774;
		3599: SAMPLE = 16'ha798;
		3600: SAMPLE = 16'ha7bd;
		3601: SAMPLE = 16'ha7e1;
		3602: SAMPLE = 16'ha806;
		3603: SAMPLE = 16'ha82a;
		3604: SAMPLE = 16'ha84f;
		3605: SAMPLE = 16'ha873;
		3606: SAMPLE = 16'ha898;
		3607: SAMPLE = 16'ha8bd;
		3608: SAMPLE = 16'ha8e2;
		3609: SAMPLE = 16'ha906;
		3610: SAMPLE = 16'ha92b;
		3611: SAMPLE = 16'ha950;
		3612: SAMPLE = 16'ha975;
		3613: SAMPLE = 16'ha99a;
		3614: SAMPLE = 16'ha9bf;
		3615: SAMPLE = 16'ha9e5;
		3616: SAMPLE = 16'haa0a;
		3617: SAMPLE = 16'haa2f;
		3618: SAMPLE = 16'haa54;
		3619: SAMPLE = 16'haa7a;
		3620: SAMPLE = 16'haa9f;
		3621: SAMPLE = 16'haac5;
		3622: SAMPLE = 16'haaea;
		3623: SAMPLE = 16'hab10;
		3624: SAMPLE = 16'hab35;
		3625: SAMPLE = 16'hab5b;
		3626: SAMPLE = 16'hab81;
		3627: SAMPLE = 16'haba7;
		3628: SAMPLE = 16'habcc;
		3629: SAMPLE = 16'habf2;
		3630: SAMPLE = 16'hac18;
		3631: SAMPLE = 16'hac3e;
		3632: SAMPLE = 16'hac64;
		3633: SAMPLE = 16'hac8a;
		3634: SAMPLE = 16'hacb1;
		3635: SAMPLE = 16'hacd7;
		3636: SAMPLE = 16'hacfd;
		3637: SAMPLE = 16'had23;
		3638: SAMPLE = 16'had4a;
		3639: SAMPLE = 16'had70;
		3640: SAMPLE = 16'had96;
		3641: SAMPLE = 16'hadbd;
		3642: SAMPLE = 16'hade3;
		3643: SAMPLE = 16'hae0a;
		3644: SAMPLE = 16'hae31;
		3645: SAMPLE = 16'hae57;
		3646: SAMPLE = 16'hae7e;
		3647: SAMPLE = 16'haea5;
		3648: SAMPLE = 16'haecc;
		3649: SAMPLE = 16'haef3;
		3650: SAMPLE = 16'haf1a;
		3651: SAMPLE = 16'haf40;
		3652: SAMPLE = 16'haf68;
		3653: SAMPLE = 16'haf8f;
		3654: SAMPLE = 16'hafb6;
		3655: SAMPLE = 16'hafdd;
		3656: SAMPLE = 16'hb004;
		3657: SAMPLE = 16'hb02b;
		3658: SAMPLE = 16'hb053;
		3659: SAMPLE = 16'hb07a;
		3660: SAMPLE = 16'hb0a1;
		3661: SAMPLE = 16'hb0c9;
		3662: SAMPLE = 16'hb0f0;
		3663: SAMPLE = 16'hb118;
		3664: SAMPLE = 16'hb140;
		3665: SAMPLE = 16'hb167;
		3666: SAMPLE = 16'hb18f;
		3667: SAMPLE = 16'hb1b7;
		3668: SAMPLE = 16'hb1de;
		3669: SAMPLE = 16'hb206;
		3670: SAMPLE = 16'hb22e;
		3671: SAMPLE = 16'hb256;
		3672: SAMPLE = 16'hb27e;
		3673: SAMPLE = 16'hb2a6;
		3674: SAMPLE = 16'hb2ce;
		3675: SAMPLE = 16'hb2f6;
		3676: SAMPLE = 16'hb31e;
		3677: SAMPLE = 16'hb347;
		3678: SAMPLE = 16'hb36f;
		3679: SAMPLE = 16'hb397;
		3680: SAMPLE = 16'hb3c0;
		3681: SAMPLE = 16'hb3e8;
		3682: SAMPLE = 16'hb410;
		3683: SAMPLE = 16'hb439;
		3684: SAMPLE = 16'hb461;
		3685: SAMPLE = 16'hb48a;
		3686: SAMPLE = 16'hb4b3;
		3687: SAMPLE = 16'hb4db;
		3688: SAMPLE = 16'hb504;
		3689: SAMPLE = 16'hb52d;
		3690: SAMPLE = 16'hb556;
		3691: SAMPLE = 16'hb57e;
		3692: SAMPLE = 16'hb5a7;
		3693: SAMPLE = 16'hb5d0;
		3694: SAMPLE = 16'hb5f9;
		3695: SAMPLE = 16'hb622;
		3696: SAMPLE = 16'hb64b;
		3697: SAMPLE = 16'hb675;
		3698: SAMPLE = 16'hb69e;
		3699: SAMPLE = 16'hb6c7;
		3700: SAMPLE = 16'hb6f0;
		3701: SAMPLE = 16'hb719;
		3702: SAMPLE = 16'hb743;
		3703: SAMPLE = 16'hb76c;
		3704: SAMPLE = 16'hb796;
		3705: SAMPLE = 16'hb7bf;
		3706: SAMPLE = 16'hb7e9;
		3707: SAMPLE = 16'hb812;
		3708: SAMPLE = 16'hb83c;
		3709: SAMPLE = 16'hb865;
		3710: SAMPLE = 16'hb88f;
		3711: SAMPLE = 16'hb8b9;
		3712: SAMPLE = 16'hb8e3;
		3713: SAMPLE = 16'hb90c;
		3714: SAMPLE = 16'hb936;
		3715: SAMPLE = 16'hb960;
		3716: SAMPLE = 16'hb98a;
		3717: SAMPLE = 16'hb9b4;
		3718: SAMPLE = 16'hb9de;
		3719: SAMPLE = 16'hba08;
		3720: SAMPLE = 16'hba32;
		3721: SAMPLE = 16'hba5c;
		3722: SAMPLE = 16'hba87;
		3723: SAMPLE = 16'hbab1;
		3724: SAMPLE = 16'hbadb;
		3725: SAMPLE = 16'hbb05;
		3726: SAMPLE = 16'hbb30;
		3727: SAMPLE = 16'hbb5a;
		3728: SAMPLE = 16'hbb85;
		3729: SAMPLE = 16'hbbaf;
		3730: SAMPLE = 16'hbbda;
		3731: SAMPLE = 16'hbc04;
		3732: SAMPLE = 16'hbc2f;
		3733: SAMPLE = 16'hbc5a;
		3734: SAMPLE = 16'hbc84;
		3735: SAMPLE = 16'hbcaf;
		3736: SAMPLE = 16'hbcda;
		3737: SAMPLE = 16'hbd05;
		3738: SAMPLE = 16'hbd2f;
		3739: SAMPLE = 16'hbd5a;
		3740: SAMPLE = 16'hbd85;
		3741: SAMPLE = 16'hbdb0;
		3742: SAMPLE = 16'hbddb;
		3743: SAMPLE = 16'hbe06;
		3744: SAMPLE = 16'hbe31;
		3745: SAMPLE = 16'hbe5d;
		3746: SAMPLE = 16'hbe88;
		3747: SAMPLE = 16'hbeb3;
		3748: SAMPLE = 16'hbede;
		3749: SAMPLE = 16'hbf09;
		3750: SAMPLE = 16'hbf35;
		3751: SAMPLE = 16'hbf60;
		3752: SAMPLE = 16'hbf8c;
		3753: SAMPLE = 16'hbfb7;
		3754: SAMPLE = 16'hbfe2;
		3755: SAMPLE = 16'hc00e;
		3756: SAMPLE = 16'hc03a;
		3757: SAMPLE = 16'hc065;
		3758: SAMPLE = 16'hc091;
		3759: SAMPLE = 16'hc0bc;
		3760: SAMPLE = 16'hc0e8;
		3761: SAMPLE = 16'hc114;
		3762: SAMPLE = 16'hc140;
		3763: SAMPLE = 16'hc16c;
		3764: SAMPLE = 16'hc197;
		3765: SAMPLE = 16'hc1c3;
		3766: SAMPLE = 16'hc1ef;
		3767: SAMPLE = 16'hc21b;
		3768: SAMPLE = 16'hc247;
		3769: SAMPLE = 16'hc273;
		3770: SAMPLE = 16'hc29f;
		3771: SAMPLE = 16'hc2cc;
		3772: SAMPLE = 16'hc2f8;
		3773: SAMPLE = 16'hc324;
		3774: SAMPLE = 16'hc350;
		3775: SAMPLE = 16'hc37c;
		3776: SAMPLE = 16'hc3a9;
		3777: SAMPLE = 16'hc3d5;
		3778: SAMPLE = 16'hc402;
		3779: SAMPLE = 16'hc42e;
		3780: SAMPLE = 16'hc45a;
		3781: SAMPLE = 16'hc487;
		3782: SAMPLE = 16'hc4b3;
		3783: SAMPLE = 16'hc4e0;
		3784: SAMPLE = 16'hc50d;
		3785: SAMPLE = 16'hc539;
		3786: SAMPLE = 16'hc566;
		3787: SAMPLE = 16'hc593;
		3788: SAMPLE = 16'hc5bf;
		3789: SAMPLE = 16'hc5ec;
		3790: SAMPLE = 16'hc619;
		3791: SAMPLE = 16'hc646;
		3792: SAMPLE = 16'hc673;
		3793: SAMPLE = 16'hc6a0;
		3794: SAMPLE = 16'hc6cd;
		3795: SAMPLE = 16'hc6f9;
		3796: SAMPLE = 16'hc727;
		3797: SAMPLE = 16'hc754;
		3798: SAMPLE = 16'hc781;
		3799: SAMPLE = 16'hc7ae;
		3800: SAMPLE = 16'hc7db;
		3801: SAMPLE = 16'hc808;
		3802: SAMPLE = 16'hc835;
		3803: SAMPLE = 16'hc863;
		3804: SAMPLE = 16'hc890;
		3805: SAMPLE = 16'hc8bd;
		3806: SAMPLE = 16'hc8eb;
		3807: SAMPLE = 16'hc918;
		3808: SAMPLE = 16'hc945;
		3809: SAMPLE = 16'hc973;
		3810: SAMPLE = 16'hc9a0;
		3811: SAMPLE = 16'hc9ce;
		3812: SAMPLE = 16'hc9fb;
		3813: SAMPLE = 16'hca29;
		3814: SAMPLE = 16'hca57;
		3815: SAMPLE = 16'hca84;
		3816: SAMPLE = 16'hcab2;
		3817: SAMPLE = 16'hcae0;
		3818: SAMPLE = 16'hcb0d;
		3819: SAMPLE = 16'hcb3b;
		3820: SAMPLE = 16'hcb69;
		3821: SAMPLE = 16'hcb97;
		3822: SAMPLE = 16'hcbc5;
		3823: SAMPLE = 16'hcbf3;
		3824: SAMPLE = 16'hcc21;
		3825: SAMPLE = 16'hcc4f;
		3826: SAMPLE = 16'hcc7d;
		3827: SAMPLE = 16'hccab;
		3828: SAMPLE = 16'hccd9;
		3829: SAMPLE = 16'hcd07;
		3830: SAMPLE = 16'hcd35;
		3831: SAMPLE = 16'hcd63;
		3832: SAMPLE = 16'hcd91;
		3833: SAMPLE = 16'hcdbf;
		3834: SAMPLE = 16'hcdee;
		3835: SAMPLE = 16'hce1c;
		3836: SAMPLE = 16'hce4a;
		3837: SAMPLE = 16'hce79;
		3838: SAMPLE = 16'hcea7;
		3839: SAMPLE = 16'hced5;
		3840: SAMPLE = 16'hcf04;
		3841: SAMPLE = 16'hcf32;
		3842: SAMPLE = 16'hcf61;
		3843: SAMPLE = 16'hcf8f;
		3844: SAMPLE = 16'hcfbe;
		3845: SAMPLE = 16'hcfec;
		3846: SAMPLE = 16'hd01b;
		3847: SAMPLE = 16'hd04a;
		3848: SAMPLE = 16'hd078;
		3849: SAMPLE = 16'hd0a7;
		3850: SAMPLE = 16'hd0d6;
		3851: SAMPLE = 16'hd104;
		3852: SAMPLE = 16'hd133;
		3853: SAMPLE = 16'hd162;
		3854: SAMPLE = 16'hd191;
		3855: SAMPLE = 16'hd1c0;
		3856: SAMPLE = 16'hd1ee;
		3857: SAMPLE = 16'hd21d;
		3858: SAMPLE = 16'hd24c;
		3859: SAMPLE = 16'hd27b;
		3860: SAMPLE = 16'hd2aa;
		3861: SAMPLE = 16'hd2d9;
		3862: SAMPLE = 16'hd308;
		3863: SAMPLE = 16'hd337;
		3864: SAMPLE = 16'hd367;
		3865: SAMPLE = 16'hd396;
		3866: SAMPLE = 16'hd3c5;
		3867: SAMPLE = 16'hd3f4;
		3868: SAMPLE = 16'hd423;
		3869: SAMPLE = 16'hd452;
		3870: SAMPLE = 16'hd482;
		3871: SAMPLE = 16'hd4b1;
		3872: SAMPLE = 16'hd4e0;
		3873: SAMPLE = 16'hd510;
		3874: SAMPLE = 16'hd53f;
		3875: SAMPLE = 16'hd56e;
		3876: SAMPLE = 16'hd59e;
		3877: SAMPLE = 16'hd5cd;
		3878: SAMPLE = 16'hd5fd;
		3879: SAMPLE = 16'hd62c;
		3880: SAMPLE = 16'hd65c;
		3881: SAMPLE = 16'hd68b;
		3882: SAMPLE = 16'hd6bb;
		3883: SAMPLE = 16'hd6ea;
		3884: SAMPLE = 16'hd71a;
		3885: SAMPLE = 16'hd74a;
		3886: SAMPLE = 16'hd779;
		3887: SAMPLE = 16'hd7a9;
		3888: SAMPLE = 16'hd7d9;
		3889: SAMPLE = 16'hd809;
		3890: SAMPLE = 16'hd838;
		3891: SAMPLE = 16'hd868;
		3892: SAMPLE = 16'hd898;
		3893: SAMPLE = 16'hd8c8;
		3894: SAMPLE = 16'hd8f8;
		3895: SAMPLE = 16'hd927;
		3896: SAMPLE = 16'hd957;
		3897: SAMPLE = 16'hd987;
		3898: SAMPLE = 16'hd9b7;
		3899: SAMPLE = 16'hd9e7;
		3900: SAMPLE = 16'hda17;
		3901: SAMPLE = 16'hda47;
		3902: SAMPLE = 16'hda77;
		3903: SAMPLE = 16'hdaa7;
		3904: SAMPLE = 16'hdad7;
		3905: SAMPLE = 16'hdb08;
		3906: SAMPLE = 16'hdb38;
		3907: SAMPLE = 16'hdb68;
		3908: SAMPLE = 16'hdb98;
		3909: SAMPLE = 16'hdbc8;
		3910: SAMPLE = 16'hdbf8;
		3911: SAMPLE = 16'hdc29;
		3912: SAMPLE = 16'hdc59;
		3913: SAMPLE = 16'hdc89;
		3914: SAMPLE = 16'hdcba;
		3915: SAMPLE = 16'hdcea;
		3916: SAMPLE = 16'hdd1a;
		3917: SAMPLE = 16'hdd4b;
		3918: SAMPLE = 16'hdd7b;
		3919: SAMPLE = 16'hddab;
		3920: SAMPLE = 16'hdddc;
		3921: SAMPLE = 16'hde0c;
		3922: SAMPLE = 16'hde3d;
		3923: SAMPLE = 16'hde6d;
		3924: SAMPLE = 16'hde9e;
		3925: SAMPLE = 16'hdece;
		3926: SAMPLE = 16'hdeff;
		3927: SAMPLE = 16'hdf2f;
		3928: SAMPLE = 16'hdf60;
		3929: SAMPLE = 16'hdf91;
		3930: SAMPLE = 16'hdfc1;
		3931: SAMPLE = 16'hdff2;
		3932: SAMPLE = 16'he023;
		3933: SAMPLE = 16'he053;
		3934: SAMPLE = 16'he084;
		3935: SAMPLE = 16'he0b5;
		3936: SAMPLE = 16'he0e6;
		3937: SAMPLE = 16'he116;
		3938: SAMPLE = 16'he147;
		3939: SAMPLE = 16'he178;
		3940: SAMPLE = 16'he1a9;
		3941: SAMPLE = 16'he1da;
		3942: SAMPLE = 16'he20a;
		3943: SAMPLE = 16'he23b;
		3944: SAMPLE = 16'he26c;
		3945: SAMPLE = 16'he29d;
		3946: SAMPLE = 16'he2ce;
		3947: SAMPLE = 16'he2ff;
		3948: SAMPLE = 16'he330;
		3949: SAMPLE = 16'he361;
		3950: SAMPLE = 16'he392;
		3951: SAMPLE = 16'he3c3;
		3952: SAMPLE = 16'he3f4;
		3953: SAMPLE = 16'he425;
		3954: SAMPLE = 16'he456;
		3955: SAMPLE = 16'he487;
		3956: SAMPLE = 16'he4b8;
		3957: SAMPLE = 16'he4e9;
		3958: SAMPLE = 16'he51b;
		3959: SAMPLE = 16'he54c;
		3960: SAMPLE = 16'he57d;
		3961: SAMPLE = 16'he5ae;
		3962: SAMPLE = 16'he5df;
		3963: SAMPLE = 16'he610;
		3964: SAMPLE = 16'he642;
		3965: SAMPLE = 16'he673;
		3966: SAMPLE = 16'he6a4;
		3967: SAMPLE = 16'he6d5;
		3968: SAMPLE = 16'he707;
		3969: SAMPLE = 16'he738;
		3970: SAMPLE = 16'he769;
		3971: SAMPLE = 16'he79b;
		3972: SAMPLE = 16'he7cc;
		3973: SAMPLE = 16'he7fd;
		3974: SAMPLE = 16'he82f;
		3975: SAMPLE = 16'he860;
		3976: SAMPLE = 16'he892;
		3977: SAMPLE = 16'he8c3;
		3978: SAMPLE = 16'he8f5;
		3979: SAMPLE = 16'he926;
		3980: SAMPLE = 16'he957;
		3981: SAMPLE = 16'he989;
		3982: SAMPLE = 16'he9ba;
		3983: SAMPLE = 16'he9ec;
		3984: SAMPLE = 16'hea1d;
		3985: SAMPLE = 16'hea4f;
		3986: SAMPLE = 16'hea80;
		3987: SAMPLE = 16'heab2;
		3988: SAMPLE = 16'heae4;
		3989: SAMPLE = 16'heb15;
		3990: SAMPLE = 16'heb47;
		3991: SAMPLE = 16'heb78;
		3992: SAMPLE = 16'hebaa;
		3993: SAMPLE = 16'hebdc;
		3994: SAMPLE = 16'hec0d;
		3995: SAMPLE = 16'hec3f;
		3996: SAMPLE = 16'hec71;
		3997: SAMPLE = 16'heca2;
		3998: SAMPLE = 16'hecd4;
		3999: SAMPLE = 16'hed06;
		4000: SAMPLE = 16'hed37;
		4001: SAMPLE = 16'hed69;
		4002: SAMPLE = 16'hed9b;
		4003: SAMPLE = 16'hedcd;
		4004: SAMPLE = 16'hedfe;
		4005: SAMPLE = 16'hee30;
		4006: SAMPLE = 16'hee62;
		4007: SAMPLE = 16'hee94;
		4008: SAMPLE = 16'heec6;
		4009: SAMPLE = 16'heef7;
		4010: SAMPLE = 16'hef29;
		4011: SAMPLE = 16'hef5b;
		4012: SAMPLE = 16'hef8d;
		4013: SAMPLE = 16'hefbf;
		4014: SAMPLE = 16'heff1;
		4015: SAMPLE = 16'hf022;
		4016: SAMPLE = 16'hf054;
		4017: SAMPLE = 16'hf086;
		4018: SAMPLE = 16'hf0b8;
		4019: SAMPLE = 16'hf0ea;
		4020: SAMPLE = 16'hf11c;
		4021: SAMPLE = 16'hf14e;
		4022: SAMPLE = 16'hf180;
		4023: SAMPLE = 16'hf1b2;
		4024: SAMPLE = 16'hf1e4;
		4025: SAMPLE = 16'hf216;
		4026: SAMPLE = 16'hf248;
		4027: SAMPLE = 16'hf27a;
		4028: SAMPLE = 16'hf2ac;
		4029: SAMPLE = 16'hf2de;
		4030: SAMPLE = 16'hf310;
		4031: SAMPLE = 16'hf342;
		4032: SAMPLE = 16'hf374;
		4033: SAMPLE = 16'hf3a6;
		4034: SAMPLE = 16'hf3d8;
		4035: SAMPLE = 16'hf40a;
		4036: SAMPLE = 16'hf43c;
		4037: SAMPLE = 16'hf46e;
		4038: SAMPLE = 16'hf4a0;
		4039: SAMPLE = 16'hf4d2;
		4040: SAMPLE = 16'hf504;
		4041: SAMPLE = 16'hf536;
		4042: SAMPLE = 16'hf568;
		4043: SAMPLE = 16'hf59a;
		4044: SAMPLE = 16'hf5cc;
		4045: SAMPLE = 16'hf5ff;
		4046: SAMPLE = 16'hf631;
		4047: SAMPLE = 16'hf663;
		4048: SAMPLE = 16'hf695;
		4049: SAMPLE = 16'hf6c7;
		4050: SAMPLE = 16'hf6f9;
		4051: SAMPLE = 16'hf72b;
		4052: SAMPLE = 16'hf75d;
		4053: SAMPLE = 16'hf790;
		4054: SAMPLE = 16'hf7c2;
		4055: SAMPLE = 16'hf7f4;
		4056: SAMPLE = 16'hf826;
		4057: SAMPLE = 16'hf858;
		4058: SAMPLE = 16'hf88a;
		4059: SAMPLE = 16'hf8bd;
		4060: SAMPLE = 16'hf8ef;
		4061: SAMPLE = 16'hf921;
		4062: SAMPLE = 16'hf953;
		4063: SAMPLE = 16'hf985;
		4064: SAMPLE = 16'hf9b8;
		4065: SAMPLE = 16'hf9ea;
		4066: SAMPLE = 16'hfa1c;
		4067: SAMPLE = 16'hfa4e;
		4068: SAMPLE = 16'hfa80;
		4069: SAMPLE = 16'hfab3;
		4070: SAMPLE = 16'hfae5;
		4071: SAMPLE = 16'hfb17;
		4072: SAMPLE = 16'hfb49;
		4073: SAMPLE = 16'hfb7c;
		4074: SAMPLE = 16'hfbae;
		4075: SAMPLE = 16'hfbe0;
		4076: SAMPLE = 16'hfc12;
		4077: SAMPLE = 16'hfc45;
		4078: SAMPLE = 16'hfc77;
		4079: SAMPLE = 16'hfca9;
		4080: SAMPLE = 16'hfcdb;
		4081: SAMPLE = 16'hfd0e;
		4082: SAMPLE = 16'hfd40;
		4083: SAMPLE = 16'hfd72;
		4084: SAMPLE = 16'hfda4;
		4085: SAMPLE = 16'hfdd7;
		4086: SAMPLE = 16'hfe09;
		4087: SAMPLE = 16'hfe3b;
		4088: SAMPLE = 16'hfe6d;
		4089: SAMPLE = 16'hfea0;
		4090: SAMPLE = 16'hfed2;
		4091: SAMPLE = 16'hff04;
		4092: SAMPLE = 16'hff36;
		4093: SAMPLE = 16'hff69;
		4094: SAMPLE = 16'hff9b;
		4095: SAMPLE = 16'hffcd;
				4096: SAMPLE = 16'h0;
		4097: SAMPLE = 16'h0;
		4098: SAMPLE = 16'h0;
		4099: SAMPLE = 16'h0;
		4100: SAMPLE = 16'h0;
		4101: SAMPLE = 16'h0;
		4102: SAMPLE = 16'h0;
		4103: SAMPLE = 16'h1;
		4104: SAMPLE = 16'h1;
		4105: SAMPLE = 16'h2;
		4106: SAMPLE = 16'h3;
		4107: SAMPLE = 16'h4;
		4108: SAMPLE = 16'h5;
		4109: SAMPLE = 16'h7;
		4110: SAMPLE = 16'h8;
		4111: SAMPLE = 16'ha;
		4112: SAMPLE = 16'hd;
		4113: SAMPLE = 16'hf;
		4114: SAMPLE = 16'h12;
		4115: SAMPLE = 16'h16;
		4116: SAMPLE = 16'h19;
		4117: SAMPLE = 16'h1d;
		4118: SAMPLE = 16'h22;
		4119: SAMPLE = 16'h26;
		4120: SAMPLE = 16'h2b;
		4121: SAMPLE = 16'h31;
		4122: SAMPLE = 16'h37;
		4123: SAMPLE = 16'h3d;
		4124: SAMPLE = 16'h44;
		4125: SAMPLE = 16'h4b;
		4126: SAMPLE = 16'h53;
		4127: SAMPLE = 16'h5c;
		4128: SAMPLE = 16'h64;
		4129: SAMPLE = 16'h6e;
		4130: SAMPLE = 16'h77;
		4131: SAMPLE = 16'h82;
		4132: SAMPLE = 16'h8c;
		4133: SAMPLE = 16'h98;
		4134: SAMPLE = 16'ha3;
		4135: SAMPLE = 16'hb0;
		4136: SAMPLE = 16'hbc;
		4137: SAMPLE = 16'hca;
		4138: SAMPLE = 16'hd8;
		4139: SAMPLE = 16'he6;
		4140: SAMPLE = 16'hf5;
		4141: SAMPLE = 16'h105;
		4142: SAMPLE = 16'h115;
		4143: SAMPLE = 16'h125;
		4144: SAMPLE = 16'h136;
		4145: SAMPLE = 16'h148;
		4146: SAMPLE = 16'h15a;
		4147: SAMPLE = 16'h16c;
		4148: SAMPLE = 16'h17f;
		4149: SAMPLE = 16'h193;
		4150: SAMPLE = 16'h1a7;
		4151: SAMPLE = 16'h1bc;
		4152: SAMPLE = 16'h1d1;
		4153: SAMPLE = 16'h1e6;
		4154: SAMPLE = 16'h1fc;
		4155: SAMPLE = 16'h212;
		4156: SAMPLE = 16'h229;
		4157: SAMPLE = 16'h240;
		4158: SAMPLE = 16'h258;
		4159: SAMPLE = 16'h26f;
		4160: SAMPLE = 16'h288;
		4161: SAMPLE = 16'h2a0;
		4162: SAMPLE = 16'h2b9;
		4163: SAMPLE = 16'h2d3;
		4164: SAMPLE = 16'h2ec;
		4165: SAMPLE = 16'h306;
		4166: SAMPLE = 16'h320;
		4167: SAMPLE = 16'h33b;
		4168: SAMPLE = 16'h356;
		4169: SAMPLE = 16'h371;
		4170: SAMPLE = 16'h38c;
		4171: SAMPLE = 16'h3a7;
		4172: SAMPLE = 16'h3c2;
		4173: SAMPLE = 16'h3de;
		4174: SAMPLE = 16'h3fa;
		4175: SAMPLE = 16'h416;
		4176: SAMPLE = 16'h432;
		4177: SAMPLE = 16'h44e;
		4178: SAMPLE = 16'h46a;
		4179: SAMPLE = 16'h486;
		4180: SAMPLE = 16'h4a2;
		4181: SAMPLE = 16'h4be;
		4182: SAMPLE = 16'h4da;
		4183: SAMPLE = 16'h4f6;
		4184: SAMPLE = 16'h512;
		4185: SAMPLE = 16'h52e;
		4186: SAMPLE = 16'h54a;
		4187: SAMPLE = 16'h566;
		4188: SAMPLE = 16'h581;
		4189: SAMPLE = 16'h59c;
		4190: SAMPLE = 16'h5b8;
		4191: SAMPLE = 16'h5d3;
		4192: SAMPLE = 16'h5ed;
		4193: SAMPLE = 16'h608;
		4194: SAMPLE = 16'h622;
		4195: SAMPLE = 16'h63c;
		4196: SAMPLE = 16'h656;
		4197: SAMPLE = 16'h66f;
		4198: SAMPLE = 16'h688;
		4199: SAMPLE = 16'h6a1;
		4200: SAMPLE = 16'h6b9;
		4201: SAMPLE = 16'h6d1;
		4202: SAMPLE = 16'h6e9;
		4203: SAMPLE = 16'h700;
		4204: SAMPLE = 16'h717;
		4205: SAMPLE = 16'h72e;
		4206: SAMPLE = 16'h744;
		4207: SAMPLE = 16'h759;
		4208: SAMPLE = 16'h76e;
		4209: SAMPLE = 16'h783;
		4210: SAMPLE = 16'h797;
		4211: SAMPLE = 16'h7ab;
		4212: SAMPLE = 16'h7be;
		4213: SAMPLE = 16'h7d0;
		4214: SAMPLE = 16'h7e3;
		4215: SAMPLE = 16'h7f4;
		4216: SAMPLE = 16'h805;
		4217: SAMPLE = 16'h816;
		4218: SAMPLE = 16'h826;
		4219: SAMPLE = 16'h836;
		4220: SAMPLE = 16'h845;
		4221: SAMPLE = 16'h853;
		4222: SAMPLE = 16'h861;
		4223: SAMPLE = 16'h86f;
		4224: SAMPLE = 16'h87c;
		4225: SAMPLE = 16'h888;
		4226: SAMPLE = 16'h894;
		4227: SAMPLE = 16'h89f;
		4228: SAMPLE = 16'h8aa;
		4229: SAMPLE = 16'h8b4;
		4230: SAMPLE = 16'h8be;
		4231: SAMPLE = 16'h8c8;
		4232: SAMPLE = 16'h8d0;
		4233: SAMPLE = 16'h8d9;
		4234: SAMPLE = 16'h8e1;
		4235: SAMPLE = 16'h8e8;
		4236: SAMPLE = 16'h8ef;
		4237: SAMPLE = 16'h8f5;
		4238: SAMPLE = 16'h8fb;
		4239: SAMPLE = 16'h901;
		4240: SAMPLE = 16'h906;
		4241: SAMPLE = 16'h90b;
		4242: SAMPLE = 16'h90f;
		4243: SAMPLE = 16'h913;
		4244: SAMPLE = 16'h917;
		4245: SAMPLE = 16'h91a;
		4246: SAMPLE = 16'h91d;
		4247: SAMPLE = 16'h91f;
		4248: SAMPLE = 16'h922;
		4249: SAMPLE = 16'h924;
		4250: SAMPLE = 16'h925;
		4251: SAMPLE = 16'h927;
		4252: SAMPLE = 16'h928;
		4253: SAMPLE = 16'h929;
		4254: SAMPLE = 16'h92a;
		4255: SAMPLE = 16'h92b;
		4256: SAMPLE = 16'h92b;
		4257: SAMPLE = 16'h92c;
		4258: SAMPLE = 16'h92c;
		4259: SAMPLE = 16'h92c;
		4260: SAMPLE = 16'h92c;
		4261: SAMPLE = 16'h92c;
		4262: SAMPLE = 16'h92c;
		4263: SAMPLE = 16'h92c;
		4264: SAMPLE = 16'h92c;
		4265: SAMPLE = 16'h92b;
		4266: SAMPLE = 16'h92b;
		4267: SAMPLE = 16'h92b;
		4268: SAMPLE = 16'h92b;
		4269: SAMPLE = 16'h92c;
		4270: SAMPLE = 16'h92c;
		4271: SAMPLE = 16'h92c;
		4272: SAMPLE = 16'h92d;
		4273: SAMPLE = 16'h92e;
		4274: SAMPLE = 16'h92e;
		4275: SAMPLE = 16'h930;
		4276: SAMPLE = 16'h931;
		4277: SAMPLE = 16'h933;
		4278: SAMPLE = 16'h934;
		4279: SAMPLE = 16'h937;
		4280: SAMPLE = 16'h939;
		4281: SAMPLE = 16'h93c;
		4282: SAMPLE = 16'h93f;
		4283: SAMPLE = 16'h942;
		4284: SAMPLE = 16'h946;
		4285: SAMPLE = 16'h94a;
		4286: SAMPLE = 16'h94f;
		4287: SAMPLE = 16'h954;
		4288: SAMPLE = 16'h959;
		4289: SAMPLE = 16'h95f;
		4290: SAMPLE = 16'h965;
		4291: SAMPLE = 16'h96c;
		4292: SAMPLE = 16'h973;
		4293: SAMPLE = 16'h97b;
		4294: SAMPLE = 16'h983;
		4295: SAMPLE = 16'h98b;
		4296: SAMPLE = 16'h994;
		4297: SAMPLE = 16'h99e;
		4298: SAMPLE = 16'h9a8;
		4299: SAMPLE = 16'h9b3;
		4300: SAMPLE = 16'h9be;
		4301: SAMPLE = 16'h9ca;
		4302: SAMPLE = 16'h9d6;
		4303: SAMPLE = 16'h9e3;
		4304: SAMPLE = 16'h9f0;
		4305: SAMPLE = 16'h9fe;
		4306: SAMPLE = 16'ha0c;
		4307: SAMPLE = 16'ha1b;
		4308: SAMPLE = 16'ha2a;
		4309: SAMPLE = 16'ha3a;
		4310: SAMPLE = 16'ha4b;
		4311: SAMPLE = 16'ha5c;
		4312: SAMPLE = 16'ha6d;
		4313: SAMPLE = 16'ha7f;
		4314: SAMPLE = 16'ha92;
		4315: SAMPLE = 16'haa5;
		4316: SAMPLE = 16'hab8;
		4317: SAMPLE = 16'hacc;
		4318: SAMPLE = 16'hae1;
		4319: SAMPLE = 16'haf6;
		4320: SAMPLE = 16'hb0b;
		4321: SAMPLE = 16'hb21;
		4322: SAMPLE = 16'hb37;
		4323: SAMPLE = 16'hb4e;
		4324: SAMPLE = 16'hb65;
		4325: SAMPLE = 16'hb7d;
		4326: SAMPLE = 16'hb95;
		4327: SAMPLE = 16'hbad;
		4328: SAMPLE = 16'hbc6;
		4329: SAMPLE = 16'hbdf;
		4330: SAMPLE = 16'hbf9;
		4331: SAMPLE = 16'hc12;
		4332: SAMPLE = 16'hc2c;
		4333: SAMPLE = 16'hc47;
		4334: SAMPLE = 16'hc61;
		4335: SAMPLE = 16'hc7c;
		4336: SAMPLE = 16'hc97;
		4337: SAMPLE = 16'hcb3;
		4338: SAMPLE = 16'hcce;
		4339: SAMPLE = 16'hcea;
		4340: SAMPLE = 16'hd06;
		4341: SAMPLE = 16'hd22;
		4342: SAMPLE = 16'hd3e;
		4343: SAMPLE = 16'hd5a;
		4344: SAMPLE = 16'hd76;
		4345: SAMPLE = 16'hd92;
		4346: SAMPLE = 16'hdaf;
		4347: SAMPLE = 16'hdcb;
		4348: SAMPLE = 16'hde7;
		4349: SAMPLE = 16'he04;
		4350: SAMPLE = 16'he20;
		4351: SAMPLE = 16'he3c;
		4352: SAMPLE = 16'he58;
		4353: SAMPLE = 16'he74;
		4354: SAMPLE = 16'he90;
		4355: SAMPLE = 16'heac;
		4356: SAMPLE = 16'hec8;
		4357: SAMPLE = 16'hee3;
		4358: SAMPLE = 16'hefe;
		4359: SAMPLE = 16'hf19;
		4360: SAMPLE = 16'hf34;
		4361: SAMPLE = 16'hf4f;
		4362: SAMPLE = 16'hf69;
		4363: SAMPLE = 16'hf83;
		4364: SAMPLE = 16'hf9d;
		4365: SAMPLE = 16'hfb6;
		4366: SAMPLE = 16'hfcf;
		4367: SAMPLE = 16'hfe8;
		4368: SAMPLE = 16'h1000;
		4369: SAMPLE = 16'h1018;
		4370: SAMPLE = 16'h102f;
		4371: SAMPLE = 16'h1046;
		4372: SAMPLE = 16'h105d;
		4373: SAMPLE = 16'h1073;
		4374: SAMPLE = 16'h1089;
		4375: SAMPLE = 16'h109e;
		4376: SAMPLE = 16'h10b3;
		4377: SAMPLE = 16'h10c7;
		4378: SAMPLE = 16'h10db;
		4379: SAMPLE = 16'h10ef;
		4380: SAMPLE = 16'h1102;
		4381: SAMPLE = 16'h1114;
		4382: SAMPLE = 16'h1126;
		4383: SAMPLE = 16'h1137;
		4384: SAMPLE = 16'h1148;
		4385: SAMPLE = 16'h1158;
		4386: SAMPLE = 16'h1168;
		4387: SAMPLE = 16'h1177;
		4388: SAMPLE = 16'h1186;
		4389: SAMPLE = 16'h1194;
		4390: SAMPLE = 16'h11a1;
		4391: SAMPLE = 16'h11ae;
		4392: SAMPLE = 16'h11bb;
		4393: SAMPLE = 16'h11c7;
		4394: SAMPLE = 16'h11d2;
		4395: SAMPLE = 16'h11dd;
		4396: SAMPLE = 16'h11e7;
		4397: SAMPLE = 16'h11f1;
		4398: SAMPLE = 16'h11fa;
		4399: SAMPLE = 16'h1203;
		4400: SAMPLE = 16'h120b;
		4401: SAMPLE = 16'h1213;
		4402: SAMPLE = 16'h121b;
		4403: SAMPLE = 16'h1221;
		4404: SAMPLE = 16'h1228;
		4405: SAMPLE = 16'h122e;
		4406: SAMPLE = 16'h1233;
		4407: SAMPLE = 16'h1238;
		4408: SAMPLE = 16'h123d;
		4409: SAMPLE = 16'h1241;
		4410: SAMPLE = 16'h1245;
		4411: SAMPLE = 16'h1248;
		4412: SAMPLE = 16'h124b;
		4413: SAMPLE = 16'h124e;
		4414: SAMPLE = 16'h1250;
		4415: SAMPLE = 16'h1252;
		4416: SAMPLE = 16'h1254;
		4417: SAMPLE = 16'h1256;
		4418: SAMPLE = 16'h1257;
		4419: SAMPLE = 16'h1258;
		4420: SAMPLE = 16'h1259;
		4421: SAMPLE = 16'h1259;
		4422: SAMPLE = 16'h125a;
		4423: SAMPLE = 16'h125a;
		4424: SAMPLE = 16'h125a;
		4425: SAMPLE = 16'h125a;
		4426: SAMPLE = 16'h1259;
		4427: SAMPLE = 16'h1259;
		4428: SAMPLE = 16'h1259;
		4429: SAMPLE = 16'h1258;
		4430: SAMPLE = 16'h1258;
		4431: SAMPLE = 16'h1257;
		4432: SAMPLE = 16'h1257;
		4433: SAMPLE = 16'h1256;
		4434: SAMPLE = 16'h1256;
		4435: SAMPLE = 16'h1256;
		4436: SAMPLE = 16'h1256;
		4437: SAMPLE = 16'h1255;
		4438: SAMPLE = 16'h1255;
		4439: SAMPLE = 16'h1256;
		4440: SAMPLE = 16'h1256;
		4441: SAMPLE = 16'h1256;
		4442: SAMPLE = 16'h1257;
		4443: SAMPLE = 16'h1258;
		4444: SAMPLE = 16'h1259;
		4445: SAMPLE = 16'h125b;
		4446: SAMPLE = 16'h125d;
		4447: SAMPLE = 16'h125f;
		4448: SAMPLE = 16'h1261;
		4449: SAMPLE = 16'h1264;
		4450: SAMPLE = 16'h1267;
		4451: SAMPLE = 16'h126a;
		4452: SAMPLE = 16'h126e;
		4453: SAMPLE = 16'h1272;
		4454: SAMPLE = 16'h1277;
		4455: SAMPLE = 16'h127c;
		4456: SAMPLE = 16'h1282;
		4457: SAMPLE = 16'h1288;
		4458: SAMPLE = 16'h128e;
		4459: SAMPLE = 16'h1295;
		4460: SAMPLE = 16'h129c;
		4461: SAMPLE = 16'h12a4;
		4462: SAMPLE = 16'h12ac;
		4463: SAMPLE = 16'h12b5;
		4464: SAMPLE = 16'h12bf;
		4465: SAMPLE = 16'h12c9;
		4466: SAMPLE = 16'h12d3;
		4467: SAMPLE = 16'h12de;
		4468: SAMPLE = 16'h12e9;
		4469: SAMPLE = 16'h12f5;
		4470: SAMPLE = 16'h1302;
		4471: SAMPLE = 16'h130f;
		4472: SAMPLE = 16'h131d;
		4473: SAMPLE = 16'h132b;
		4474: SAMPLE = 16'h133a;
		4475: SAMPLE = 16'h1349;
		4476: SAMPLE = 16'h1359;
		4477: SAMPLE = 16'h136a;
		4478: SAMPLE = 16'h137b;
		4479: SAMPLE = 16'h138c;
		4480: SAMPLE = 16'h139e;
		4481: SAMPLE = 16'h13b1;
		4482: SAMPLE = 16'h13c4;
		4483: SAMPLE = 16'h13d7;
		4484: SAMPLE = 16'h13ec;
		4485: SAMPLE = 16'h1400;
		4486: SAMPLE = 16'h1415;
		4487: SAMPLE = 16'h142b;
		4488: SAMPLE = 16'h1441;
		4489: SAMPLE = 16'h1457;
		4490: SAMPLE = 16'h146e;
		4491: SAMPLE = 16'h1486;
		4492: SAMPLE = 16'h149e;
		4493: SAMPLE = 16'h14b6;
		4494: SAMPLE = 16'h14cf;
		4495: SAMPLE = 16'h14e8;
		4496: SAMPLE = 16'h1501;
		4497: SAMPLE = 16'h151b;
		4498: SAMPLE = 16'h1535;
		4499: SAMPLE = 16'h154f;
		4500: SAMPLE = 16'h156a;
		4501: SAMPLE = 16'h1585;
		4502: SAMPLE = 16'h15a0;
		4503: SAMPLE = 16'h15bb;
		4504: SAMPLE = 16'h15d7;
		4505: SAMPLE = 16'h15f3;
		4506: SAMPLE = 16'h160f;
		4507: SAMPLE = 16'h162b;
		4508: SAMPLE = 16'h1648;
		4509: SAMPLE = 16'h1664;
		4510: SAMPLE = 16'h1681;
		4511: SAMPLE = 16'h169e;
		4512: SAMPLE = 16'h16ba;
		4513: SAMPLE = 16'h16d7;
		4514: SAMPLE = 16'h16f4;
		4515: SAMPLE = 16'h1711;
		4516: SAMPLE = 16'h172e;
		4517: SAMPLE = 16'h174b;
		4518: SAMPLE = 16'h1767;
		4519: SAMPLE = 16'h1784;
		4520: SAMPLE = 16'h17a1;
		4521: SAMPLE = 16'h17bd;
		4522: SAMPLE = 16'h17d9;
		4523: SAMPLE = 16'h17f5;
		4524: SAMPLE = 16'h1811;
		4525: SAMPLE = 16'h182d;
		4526: SAMPLE = 16'h1849;
		4527: SAMPLE = 16'h1864;
		4528: SAMPLE = 16'h187f;
		4529: SAMPLE = 16'h189a;
		4530: SAMPLE = 16'h18b4;
		4531: SAMPLE = 16'h18ce;
		4532: SAMPLE = 16'h18e8;
		4533: SAMPLE = 16'h1901;
		4534: SAMPLE = 16'h191b;
		4535: SAMPLE = 16'h1933;
		4536: SAMPLE = 16'h194c;
		4537: SAMPLE = 16'h1964;
		4538: SAMPLE = 16'h197b;
		4539: SAMPLE = 16'h1992;
		4540: SAMPLE = 16'h19a9;
		4541: SAMPLE = 16'h19bf;
		4542: SAMPLE = 16'h19d4;
		4543: SAMPLE = 16'h19ea;
		4544: SAMPLE = 16'h19fe;
		4545: SAMPLE = 16'h1a13;
		4546: SAMPLE = 16'h1a26;
		4547: SAMPLE = 16'h1a39;
		4548: SAMPLE = 16'h1a4c;
		4549: SAMPLE = 16'h1a5e;
		4550: SAMPLE = 16'h1a70;
		4551: SAMPLE = 16'h1a81;
		4552: SAMPLE = 16'h1a91;
		4553: SAMPLE = 16'h1aa1;
		4554: SAMPLE = 16'h1ab0;
		4555: SAMPLE = 16'h1abf;
		4556: SAMPLE = 16'h1acd;
		4557: SAMPLE = 16'h1adb;
		4558: SAMPLE = 16'h1ae8;
		4559: SAMPLE = 16'h1af4;
		4560: SAMPLE = 16'h1b00;
		4561: SAMPLE = 16'h1b0c;
		4562: SAMPLE = 16'h1b16;
		4563: SAMPLE = 16'h1b21;
		4564: SAMPLE = 16'h1b2b;
		4565: SAMPLE = 16'h1b34;
		4566: SAMPLE = 16'h1b3c;
		4567: SAMPLE = 16'h1b45;
		4568: SAMPLE = 16'h1b4c;
		4569: SAMPLE = 16'h1b53;
		4570: SAMPLE = 16'h1b5a;
		4571: SAMPLE = 16'h1b60;
		4572: SAMPLE = 16'h1b66;
		4573: SAMPLE = 16'h1b6b;
		4574: SAMPLE = 16'h1b70;
		4575: SAMPLE = 16'h1b74;
		4576: SAMPLE = 16'h1b78;
		4577: SAMPLE = 16'h1b7b;
		4578: SAMPLE = 16'h1b7e;
		4579: SAMPLE = 16'h1b81;
		4580: SAMPLE = 16'h1b83;
		4581: SAMPLE = 16'h1b85;
		4582: SAMPLE = 16'h1b87;
		4583: SAMPLE = 16'h1b88;
		4584: SAMPLE = 16'h1b89;
		4585: SAMPLE = 16'h1b8a;
		4586: SAMPLE = 16'h1b8b;
		4587: SAMPLE = 16'h1b8b;
		4588: SAMPLE = 16'h1b8b;
		4589: SAMPLE = 16'h1b8b;
		4590: SAMPLE = 16'h1b8a;
		4591: SAMPLE = 16'h1b8a;
		4592: SAMPLE = 16'h1b89;
		4593: SAMPLE = 16'h1b88;
		4594: SAMPLE = 16'h1b87;
		4595: SAMPLE = 16'h1b86;
		4596: SAMPLE = 16'h1b85;
		4597: SAMPLE = 16'h1b84;
		4598: SAMPLE = 16'h1b83;
		4599: SAMPLE = 16'h1b82;
		4600: SAMPLE = 16'h1b81;
		4601: SAMPLE = 16'h1b80;
		4602: SAMPLE = 16'h1b7f;
		4603: SAMPLE = 16'h1b7e;
		4604: SAMPLE = 16'h1b7d;
		4605: SAMPLE = 16'h1b7d;
		4606: SAMPLE = 16'h1b7c;
		4607: SAMPLE = 16'h1b7c;
		4608: SAMPLE = 16'h1b7c;
		4609: SAMPLE = 16'h1b7c;
		4610: SAMPLE = 16'h1b7c;
		4611: SAMPLE = 16'h1b7d;
		4612: SAMPLE = 16'h1b7e;
		4613: SAMPLE = 16'h1b7f;
		4614: SAMPLE = 16'h1b80;
		4615: SAMPLE = 16'h1b82;
		4616: SAMPLE = 16'h1b84;
		4617: SAMPLE = 16'h1b87;
		4618: SAMPLE = 16'h1b8a;
		4619: SAMPLE = 16'h1b8d;
		4620: SAMPLE = 16'h1b91;
		4621: SAMPLE = 16'h1b95;
		4622: SAMPLE = 16'h1b99;
		4623: SAMPLE = 16'h1b9e;
		4624: SAMPLE = 16'h1ba4;
		4625: SAMPLE = 16'h1baa;
		4626: SAMPLE = 16'h1bb0;
		4627: SAMPLE = 16'h1bb7;
		4628: SAMPLE = 16'h1bbf;
		4629: SAMPLE = 16'h1bc6;
		4630: SAMPLE = 16'h1bcf;
		4631: SAMPLE = 16'h1bd8;
		4632: SAMPLE = 16'h1be2;
		4633: SAMPLE = 16'h1bec;
		4634: SAMPLE = 16'h1bf7;
		4635: SAMPLE = 16'h1c02;
		4636: SAMPLE = 16'h1c0e;
		4637: SAMPLE = 16'h1c1a;
		4638: SAMPLE = 16'h1c27;
		4639: SAMPLE = 16'h1c35;
		4640: SAMPLE = 16'h1c43;
		4641: SAMPLE = 16'h1c51;
		4642: SAMPLE = 16'h1c61;
		4643: SAMPLE = 16'h1c71;
		4644: SAMPLE = 16'h1c81;
		4645: SAMPLE = 16'h1c92;
		4646: SAMPLE = 16'h1ca4;
		4647: SAMPLE = 16'h1cb6;
		4648: SAMPLE = 16'h1cc8;
		4649: SAMPLE = 16'h1cdc;
		4650: SAMPLE = 16'h1cf0;
		4651: SAMPLE = 16'h1d04;
		4652: SAMPLE = 16'h1d19;
		4653: SAMPLE = 16'h1d2e;
		4654: SAMPLE = 16'h1d44;
		4655: SAMPLE = 16'h1d5a;
		4656: SAMPLE = 16'h1d71;
		4657: SAMPLE = 16'h1d89;
		4658: SAMPLE = 16'h1da0;
		4659: SAMPLE = 16'h1db9;
		4660: SAMPLE = 16'h1dd1;
		4661: SAMPLE = 16'h1dea;
		4662: SAMPLE = 16'h1e04;
		4663: SAMPLE = 16'h1e1e;
		4664: SAMPLE = 16'h1e38;
		4665: SAMPLE = 16'h1e53;
		4666: SAMPLE = 16'h1e6e;
		4667: SAMPLE = 16'h1e89;
		4668: SAMPLE = 16'h1ea4;
		4669: SAMPLE = 16'h1ec0;
		4670: SAMPLE = 16'h1edc;
		4671: SAMPLE = 16'h1ef9;
		4672: SAMPLE = 16'h1f15;
		4673: SAMPLE = 16'h1f32;
		4674: SAMPLE = 16'h1f4f;
		4675: SAMPLE = 16'h1f6c;
		4676: SAMPLE = 16'h1f89;
		4677: SAMPLE = 16'h1fa7;
		4678: SAMPLE = 16'h1fc4;
		4679: SAMPLE = 16'h1fe2;
		4680: SAMPLE = 16'h2000;
		4681: SAMPLE = 16'h201d;
		4682: SAMPLE = 16'h203b;
		4683: SAMPLE = 16'h2058;
		4684: SAMPLE = 16'h2076;
		4685: SAMPLE = 16'h2094;
		4686: SAMPLE = 16'h20b1;
		4687: SAMPLE = 16'h20ce;
		4688: SAMPLE = 16'h20ec;
		4689: SAMPLE = 16'h2109;
		4690: SAMPLE = 16'h2126;
		4691: SAMPLE = 16'h2142;
		4692: SAMPLE = 16'h215f;
		4693: SAMPLE = 16'h217b;
		4694: SAMPLE = 16'h2197;
		4695: SAMPLE = 16'h21b3;
		4696: SAMPLE = 16'h21cf;
		4697: SAMPLE = 16'h21ea;
		4698: SAMPLE = 16'h2205;
		4699: SAMPLE = 16'h221f;
		4700: SAMPLE = 16'h2239;
		4701: SAMPLE = 16'h2253;
		4702: SAMPLE = 16'h226d;
		4703: SAMPLE = 16'h2285;
		4704: SAMPLE = 16'h229e;
		4705: SAMPLE = 16'h22b6;
		4706: SAMPLE = 16'h22ce;
		4707: SAMPLE = 16'h22e5;
		4708: SAMPLE = 16'h22fc;
		4709: SAMPLE = 16'h2312;
		4710: SAMPLE = 16'h2327;
		4711: SAMPLE = 16'h233d;
		4712: SAMPLE = 16'h2351;
		4713: SAMPLE = 16'h2365;
		4714: SAMPLE = 16'h2379;
		4715: SAMPLE = 16'h238c;
		4716: SAMPLE = 16'h239e;
		4717: SAMPLE = 16'h23b0;
		4718: SAMPLE = 16'h23c1;
		4719: SAMPLE = 16'h23d2;
		4720: SAMPLE = 16'h23e2;
		4721: SAMPLE = 16'h23f2;
		4722: SAMPLE = 16'h2401;
		4723: SAMPLE = 16'h240f;
		4724: SAMPLE = 16'h241d;
		4725: SAMPLE = 16'h242a;
		4726: SAMPLE = 16'h2436;
		4727: SAMPLE = 16'h2442;
		4728: SAMPLE = 16'h244e;
		4729: SAMPLE = 16'h2458;
		4730: SAMPLE = 16'h2462;
		4731: SAMPLE = 16'h246c;
		4732: SAMPLE = 16'h2475;
		4733: SAMPLE = 16'h247e;
		4734: SAMPLE = 16'h2485;
		4735: SAMPLE = 16'h248d;
		4736: SAMPLE = 16'h2494;
		4737: SAMPLE = 16'h249a;
		4738: SAMPLE = 16'h24a0;
		4739: SAMPLE = 16'h24a5;
		4740: SAMPLE = 16'h24aa;
		4741: SAMPLE = 16'h24ae;
		4742: SAMPLE = 16'h24b2;
		4743: SAMPLE = 16'h24b5;
		4744: SAMPLE = 16'h24b8;
		4745: SAMPLE = 16'h24ba;
		4746: SAMPLE = 16'h24bc;
		4747: SAMPLE = 16'h24be;
		4748: SAMPLE = 16'h24bf;
		4749: SAMPLE = 16'h24c0;
		4750: SAMPLE = 16'h24c1;
		4751: SAMPLE = 16'h24c1;
		4752: SAMPLE = 16'h24c1;
		4753: SAMPLE = 16'h24c1;
		4754: SAMPLE = 16'h24c0;
		4755: SAMPLE = 16'h24bf;
		4756: SAMPLE = 16'h24be;
		4757: SAMPLE = 16'h24bd;
		4758: SAMPLE = 16'h24bc;
		4759: SAMPLE = 16'h24ba;
		4760: SAMPLE = 16'h24b8;
		4761: SAMPLE = 16'h24b6;
		4762: SAMPLE = 16'h24b5;
		4763: SAMPLE = 16'h24b3;
		4764: SAMPLE = 16'h24b0;
		4765: SAMPLE = 16'h24ae;
		4766: SAMPLE = 16'h24ac;
		4767: SAMPLE = 16'h24aa;
		4768: SAMPLE = 16'h24a8;
		4769: SAMPLE = 16'h24a6;
		4770: SAMPLE = 16'h24a4;
		4771: SAMPLE = 16'h24a3;
		4772: SAMPLE = 16'h24a1;
		4773: SAMPLE = 16'h24a0;
		4774: SAMPLE = 16'h249e;
		4775: SAMPLE = 16'h249d;
		4776: SAMPLE = 16'h249d;
		4777: SAMPLE = 16'h249c;
		4778: SAMPLE = 16'h249c;
		4779: SAMPLE = 16'h249c;
		4780: SAMPLE = 16'h249c;
		4781: SAMPLE = 16'h249c;
		4782: SAMPLE = 16'h249d;
		4783: SAMPLE = 16'h249f;
		4784: SAMPLE = 16'h24a0;
		4785: SAMPLE = 16'h24a2;
		4786: SAMPLE = 16'h24a5;
		4787: SAMPLE = 16'h24a8;
		4788: SAMPLE = 16'h24ab;
		4789: SAMPLE = 16'h24af;
		4790: SAMPLE = 16'h24b3;
		4791: SAMPLE = 16'h24b8;
		4792: SAMPLE = 16'h24bd;
		4793: SAMPLE = 16'h24c3;
		4794: SAMPLE = 16'h24ca;
		4795: SAMPLE = 16'h24d1;
		4796: SAMPLE = 16'h24d8;
		4797: SAMPLE = 16'h24e0;
		4798: SAMPLE = 16'h24e9;
		4799: SAMPLE = 16'h24f2;
		4800: SAMPLE = 16'h24fc;
		4801: SAMPLE = 16'h2506;
		4802: SAMPLE = 16'h2511;
		4803: SAMPLE = 16'h251c;
		4804: SAMPLE = 16'h2529;
		4805: SAMPLE = 16'h2535;
		4806: SAMPLE = 16'h2543;
		4807: SAMPLE = 16'h2551;
		4808: SAMPLE = 16'h2560;
		4809: SAMPLE = 16'h256f;
		4810: SAMPLE = 16'h257f;
		4811: SAMPLE = 16'h258f;
		4812: SAMPLE = 16'h25a0;
		4813: SAMPLE = 16'h25b2;
		4814: SAMPLE = 16'h25c4;
		4815: SAMPLE = 16'h25d7;
		4816: SAMPLE = 16'h25eb;
		4817: SAMPLE = 16'h25ff;
		4818: SAMPLE = 16'h2614;
		4819: SAMPLE = 16'h2629;
		4820: SAMPLE = 16'h263f;
		4821: SAMPLE = 16'h2655;
		4822: SAMPLE = 16'h266c;
		4823: SAMPLE = 16'h2683;
		4824: SAMPLE = 16'h269b;
		4825: SAMPLE = 16'h26b4;
		4826: SAMPLE = 16'h26cc;
		4827: SAMPLE = 16'h26e6;
		4828: SAMPLE = 16'h2700;
		4829: SAMPLE = 16'h271a;
		4830: SAMPLE = 16'h2735;
		4831: SAMPLE = 16'h2750;
		4832: SAMPLE = 16'h276b;
		4833: SAMPLE = 16'h2787;
		4834: SAMPLE = 16'h27a3;
		4835: SAMPLE = 16'h27c0;
		4836: SAMPLE = 16'h27dc;
		4837: SAMPLE = 16'h27f9;
		4838: SAMPLE = 16'h2817;
		4839: SAMPLE = 16'h2834;
		4840: SAMPLE = 16'h2852;
		4841: SAMPLE = 16'h2870;
		4842: SAMPLE = 16'h288f;
		4843: SAMPLE = 16'h28ad;
		4844: SAMPLE = 16'h28cb;
		4845: SAMPLE = 16'h28ea;
		4846: SAMPLE = 16'h2909;
		4847: SAMPLE = 16'h2927;
		4848: SAMPLE = 16'h2946;
		4849: SAMPLE = 16'h2965;
		4850: SAMPLE = 16'h2984;
		4851: SAMPLE = 16'h29a3;
		4852: SAMPLE = 16'h29c1;
		4853: SAMPLE = 16'h29e0;
		4854: SAMPLE = 16'h29ff;
		4855: SAMPLE = 16'h2a1d;
		4856: SAMPLE = 16'h2a3b;
		4857: SAMPLE = 16'h2a59;
		4858: SAMPLE = 16'h2a77;
		4859: SAMPLE = 16'h2a95;
		4860: SAMPLE = 16'h2ab2;
		4861: SAMPLE = 16'h2ad0;
		4862: SAMPLE = 16'h2aec;
		4863: SAMPLE = 16'h2b09;
		4864: SAMPLE = 16'h2b25;
		4865: SAMPLE = 16'h2b41;
		4866: SAMPLE = 16'h2b5d;
		4867: SAMPLE = 16'h2b78;
		4868: SAMPLE = 16'h2b93;
		4869: SAMPLE = 16'h2bad;
		4870: SAMPLE = 16'h2bc7;
		4871: SAMPLE = 16'h2be0;
		4872: SAMPLE = 16'h2bf9;
		4873: SAMPLE = 16'h2c12;
		4874: SAMPLE = 16'h2c2a;
		4875: SAMPLE = 16'h2c41;
		4876: SAMPLE = 16'h2c58;
		4877: SAMPLE = 16'h2c6f;
		4878: SAMPLE = 16'h2c85;
		4879: SAMPLE = 16'h2c9a;
		4880: SAMPLE = 16'h2cae;
		4881: SAMPLE = 16'h2cc3;
		4882: SAMPLE = 16'h2cd6;
		4883: SAMPLE = 16'h2ce9;
		4884: SAMPLE = 16'h2cfb;
		4885: SAMPLE = 16'h2d0d;
		4886: SAMPLE = 16'h2d1e;
		4887: SAMPLE = 16'h2d2e;
		4888: SAMPLE = 16'h2d3e;
		4889: SAMPLE = 16'h2d4d;
		4890: SAMPLE = 16'h2d5b;
		4891: SAMPLE = 16'h2d69;
		4892: SAMPLE = 16'h2d76;
		4893: SAMPLE = 16'h2d83;
		4894: SAMPLE = 16'h2d8f;
		4895: SAMPLE = 16'h2d9a;
		4896: SAMPLE = 16'h2da5;
		4897: SAMPLE = 16'h2daf;
		4898: SAMPLE = 16'h2db8;
		4899: SAMPLE = 16'h2dc1;
		4900: SAMPLE = 16'h2dc9;
		4901: SAMPLE = 16'h2dd0;
		4902: SAMPLE = 16'h2dd7;
		4903: SAMPLE = 16'h2dde;
		4904: SAMPLE = 16'h2de3;
		4905: SAMPLE = 16'h2de8;
		4906: SAMPLE = 16'h2ded;
		4907: SAMPLE = 16'h2df1;
		4908: SAMPLE = 16'h2df5;
		4909: SAMPLE = 16'h2df8;
		4910: SAMPLE = 16'h2dfa;
		4911: SAMPLE = 16'h2dfc;
		4912: SAMPLE = 16'h2dfe;
		4913: SAMPLE = 16'h2dff;
		4914: SAMPLE = 16'h2e00;
		4915: SAMPLE = 16'h2e00;
		4916: SAMPLE = 16'h2e00;
		4917: SAMPLE = 16'h2dff;
		4918: SAMPLE = 16'h2dfe;
		4919: SAMPLE = 16'h2dfd;
		4920: SAMPLE = 16'h2dfc;
		4921: SAMPLE = 16'h2dfa;
		4922: SAMPLE = 16'h2df8;
		4923: SAMPLE = 16'h2df6;
		4924: SAMPLE = 16'h2df3;
		4925: SAMPLE = 16'h2df0;
		4926: SAMPLE = 16'h2ded;
		4927: SAMPLE = 16'h2dea;
		4928: SAMPLE = 16'h2de7;
		4929: SAMPLE = 16'h2de4;
		4930: SAMPLE = 16'h2de1;
		4931: SAMPLE = 16'h2ddd;
		4932: SAMPLE = 16'h2dda;
		4933: SAMPLE = 16'h2dd6;
		4934: SAMPLE = 16'h2dd3;
		4935: SAMPLE = 16'h2dcf;
		4936: SAMPLE = 16'h2dcc;
		4937: SAMPLE = 16'h2dc9;
		4938: SAMPLE = 16'h2dc5;
		4939: SAMPLE = 16'h2dc2;
		4940: SAMPLE = 16'h2dc0;
		4941: SAMPLE = 16'h2dbd;
		4942: SAMPLE = 16'h2dba;
		4943: SAMPLE = 16'h2db8;
		4944: SAMPLE = 16'h2db6;
		4945: SAMPLE = 16'h2db5;
		4946: SAMPLE = 16'h2db3;
		4947: SAMPLE = 16'h2db2;
		4948: SAMPLE = 16'h2db2;
		4949: SAMPLE = 16'h2db1;
		4950: SAMPLE = 16'h2db1;
		4951: SAMPLE = 16'h2db2;
		4952: SAMPLE = 16'h2db3;
		4953: SAMPLE = 16'h2db4;
		4954: SAMPLE = 16'h2db6;
		4955: SAMPLE = 16'h2db8;
		4956: SAMPLE = 16'h2dbb;
		4957: SAMPLE = 16'h2dbe;
		4958: SAMPLE = 16'h2dc2;
		4959: SAMPLE = 16'h2dc7;
		4960: SAMPLE = 16'h2dcc;
		4961: SAMPLE = 16'h2dd1;
		4962: SAMPLE = 16'h2dd7;
		4963: SAMPLE = 16'h2dde;
		4964: SAMPLE = 16'h2de5;
		4965: SAMPLE = 16'h2ded;
		4966: SAMPLE = 16'h2df6;
		4967: SAMPLE = 16'h2dff;
		4968: SAMPLE = 16'h2e09;
		4969: SAMPLE = 16'h2e14;
		4970: SAMPLE = 16'h2e1f;
		4971: SAMPLE = 16'h2e2b;
		4972: SAMPLE = 16'h2e37;
		4973: SAMPLE = 16'h2e45;
		4974: SAMPLE = 16'h2e53;
		4975: SAMPLE = 16'h2e61;
		4976: SAMPLE = 16'h2e70;
		4977: SAMPLE = 16'h2e80;
		4978: SAMPLE = 16'h2e91;
		4979: SAMPLE = 16'h2ea2;
		4980: SAMPLE = 16'h2eb4;
		4981: SAMPLE = 16'h2ec7;
		4982: SAMPLE = 16'h2eda;
		4983: SAMPLE = 16'h2eee;
		4984: SAMPLE = 16'h2f02;
		4985: SAMPLE = 16'h2f18;
		4986: SAMPLE = 16'h2f2d;
		4987: SAMPLE = 16'h2f44;
		4988: SAMPLE = 16'h2f5b;
		4989: SAMPLE = 16'h2f73;
		4990: SAMPLE = 16'h2f8b;
		4991: SAMPLE = 16'h2fa3;
		4992: SAMPLE = 16'h2fbd;
		4993: SAMPLE = 16'h2fd7;
		4994: SAMPLE = 16'h2ff1;
		4995: SAMPLE = 16'h300c;
		4996: SAMPLE = 16'h3027;
		4997: SAMPLE = 16'h3043;
		4998: SAMPLE = 16'h305f;
		4999: SAMPLE = 16'h307c;
		5000: SAMPLE = 16'h3099;
		5001: SAMPLE = 16'h30b7;
		5002: SAMPLE = 16'h30d4;
		5003: SAMPLE = 16'h30f3;
		5004: SAMPLE = 16'h3111;
		5005: SAMPLE = 16'h3130;
		5006: SAMPLE = 16'h314f;
		5007: SAMPLE = 16'h316e;
		5008: SAMPLE = 16'h318e;
		5009: SAMPLE = 16'h31ae;
		5010: SAMPLE = 16'h31ce;
		5011: SAMPLE = 16'h31ee;
		5012: SAMPLE = 16'h320e;
		5013: SAMPLE = 16'h322f;
		5014: SAMPLE = 16'h324f;
		5015: SAMPLE = 16'h326f;
		5016: SAMPLE = 16'h3290;
		5017: SAMPLE = 16'h32b0;
		5018: SAMPLE = 16'h32d1;
		5019: SAMPLE = 16'h32f1;
		5020: SAMPLE = 16'h3312;
		5021: SAMPLE = 16'h3332;
		5022: SAMPLE = 16'h3352;
		5023: SAMPLE = 16'h3372;
		5024: SAMPLE = 16'h3392;
		5025: SAMPLE = 16'h33b1;
		5026: SAMPLE = 16'h33d1;
		5027: SAMPLE = 16'h33f0;
		5028: SAMPLE = 16'h340e;
		5029: SAMPLE = 16'h342d;
		5030: SAMPLE = 16'h344b;
		5031: SAMPLE = 16'h3469;
		5032: SAMPLE = 16'h3486;
		5033: SAMPLE = 16'h34a3;
		5034: SAMPLE = 16'h34c0;
		5035: SAMPLE = 16'h34dc;
		5036: SAMPLE = 16'h34f8;
		5037: SAMPLE = 16'h3513;
		5038: SAMPLE = 16'h352e;
		5039: SAMPLE = 16'h3548;
		5040: SAMPLE = 16'h3562;
		5041: SAMPLE = 16'h357b;
		5042: SAMPLE = 16'h3593;
		5043: SAMPLE = 16'h35ab;
		5044: SAMPLE = 16'h35c3;
		5045: SAMPLE = 16'h35da;
		5046: SAMPLE = 16'h35f0;
		5047: SAMPLE = 16'h3605;
		5048: SAMPLE = 16'h361a;
		5049: SAMPLE = 16'h362e;
		5050: SAMPLE = 16'h3642;
		5051: SAMPLE = 16'h3655;
		5052: SAMPLE = 16'h3667;
		5053: SAMPLE = 16'h3678;
		5054: SAMPLE = 16'h3689;
		5055: SAMPLE = 16'h3699;
		5056: SAMPLE = 16'h36a8;
		5057: SAMPLE = 16'h36b7;
		5058: SAMPLE = 16'h36c5;
		5059: SAMPLE = 16'h36d2;
		5060: SAMPLE = 16'h36df;
		5061: SAMPLE = 16'h36ea;
		5062: SAMPLE = 16'h36f5;
		5063: SAMPLE = 16'h3700;
		5064: SAMPLE = 16'h3709;
		5065: SAMPLE = 16'h3712;
		5066: SAMPLE = 16'h371b;
		5067: SAMPLE = 16'h3722;
		5068: SAMPLE = 16'h3729;
		5069: SAMPLE = 16'h372f;
		5070: SAMPLE = 16'h3735;
		5071: SAMPLE = 16'h373a;
		5072: SAMPLE = 16'h373e;
		5073: SAMPLE = 16'h3742;
		5074: SAMPLE = 16'h3745;
		5075: SAMPLE = 16'h3747;
		5076: SAMPLE = 16'h3749;
		5077: SAMPLE = 16'h374b;
		5078: SAMPLE = 16'h374b;
		5079: SAMPLE = 16'h374c;
		5080: SAMPLE = 16'h374b;
		5081: SAMPLE = 16'h374b;
		5082: SAMPLE = 16'h374a;
		5083: SAMPLE = 16'h3748;
		5084: SAMPLE = 16'h3746;
		5085: SAMPLE = 16'h3743;
		5086: SAMPLE = 16'h3741;
		5087: SAMPLE = 16'h373d;
		5088: SAMPLE = 16'h373a;
		5089: SAMPLE = 16'h3736;
		5090: SAMPLE = 16'h3732;
		5091: SAMPLE = 16'h372e;
		5092: SAMPLE = 16'h3729;
		5093: SAMPLE = 16'h3724;
		5094: SAMPLE = 16'h371f;
		5095: SAMPLE = 16'h371a;
		5096: SAMPLE = 16'h3715;
		5097: SAMPLE = 16'h370f;
		5098: SAMPLE = 16'h370a;
		5099: SAMPLE = 16'h3704;
		5100: SAMPLE = 16'h36ff;
		5101: SAMPLE = 16'h36f9;
		5102: SAMPLE = 16'h36f4;
		5103: SAMPLE = 16'h36ee;
		5104: SAMPLE = 16'h36e9;
		5105: SAMPLE = 16'h36e4;
		5106: SAMPLE = 16'h36df;
		5107: SAMPLE = 16'h36da;
		5108: SAMPLE = 16'h36d5;
		5109: SAMPLE = 16'h36d1;
		5110: SAMPLE = 16'h36cd;
		5111: SAMPLE = 16'h36c9;
		5112: SAMPLE = 16'h36c5;
		5113: SAMPLE = 16'h36c2;
		5114: SAMPLE = 16'h36bf;
		5115: SAMPLE = 16'h36bd;
		5116: SAMPLE = 16'h36bb;
		5117: SAMPLE = 16'h36b9;
		5118: SAMPLE = 16'h36b8;
		5119: SAMPLE = 16'h36b7;
		5120: SAMPLE = 16'h36b7;
		5121: SAMPLE = 16'h36b7;
		5122: SAMPLE = 16'h36b8;
		5123: SAMPLE = 16'h36b9;
		5124: SAMPLE = 16'h36bb;
		5125: SAMPLE = 16'h36be;
		5126: SAMPLE = 16'h36c1;
		5127: SAMPLE = 16'h36c4;
		5128: SAMPLE = 16'h36c9;
		5129: SAMPLE = 16'h36ce;
		5130: SAMPLE = 16'h36d4;
		5131: SAMPLE = 16'h36da;
		5132: SAMPLE = 16'h36e1;
		5133: SAMPLE = 16'h36e9;
		5134: SAMPLE = 16'h36f2;
		5135: SAMPLE = 16'h36fb;
		5136: SAMPLE = 16'h3705;
		5137: SAMPLE = 16'h3710;
		5138: SAMPLE = 16'h371b;
		5139: SAMPLE = 16'h3727;
		5140: SAMPLE = 16'h3734;
		5141: SAMPLE = 16'h3742;
		5142: SAMPLE = 16'h3751;
		5143: SAMPLE = 16'h3760;
		5144: SAMPLE = 16'h3770;
		5145: SAMPLE = 16'h3781;
		5146: SAMPLE = 16'h3792;
		5147: SAMPLE = 16'h37a4;
		5148: SAMPLE = 16'h37b7;
		5149: SAMPLE = 16'h37cb;
		5150: SAMPLE = 16'h37e0;
		5151: SAMPLE = 16'h37f5;
		5152: SAMPLE = 16'h380b;
		5153: SAMPLE = 16'h3822;
		5154: SAMPLE = 16'h3839;
		5155: SAMPLE = 16'h3851;
		5156: SAMPLE = 16'h386a;
		5157: SAMPLE = 16'h3883;
		5158: SAMPLE = 16'h389d;
		5159: SAMPLE = 16'h38b8;
		5160: SAMPLE = 16'h38d3;
		5161: SAMPLE = 16'h38ef;
		5162: SAMPLE = 16'h390b;
		5163: SAMPLE = 16'h3928;
		5164: SAMPLE = 16'h3946;
		5165: SAMPLE = 16'h3964;
		5166: SAMPLE = 16'h3982;
		5167: SAMPLE = 16'h39a1;
		5168: SAMPLE = 16'h39c1;
		5169: SAMPLE = 16'h39e0;
		5170: SAMPLE = 16'h3a01;
		5171: SAMPLE = 16'h3a21;
		5172: SAMPLE = 16'h3a42;
		5173: SAMPLE = 16'h3a63;
		5174: SAMPLE = 16'h3a85;
		5175: SAMPLE = 16'h3aa7;
		5176: SAMPLE = 16'h3ac9;
		5177: SAMPLE = 16'h3aeb;
		5178: SAMPLE = 16'h3b0e;
		5179: SAMPLE = 16'h3b30;
		5180: SAMPLE = 16'h3b53;
		5181: SAMPLE = 16'h3b76;
		5182: SAMPLE = 16'h3b99;
		5183: SAMPLE = 16'h3bbc;
		5184: SAMPLE = 16'h3bdf;
		5185: SAMPLE = 16'h3c02;
		5186: SAMPLE = 16'h3c24;
		5187: SAMPLE = 16'h3c47;
		5188: SAMPLE = 16'h3c6a;
		5189: SAMPLE = 16'h3c8d;
		5190: SAMPLE = 16'h3caf;
		5191: SAMPLE = 16'h3cd1;
		5192: SAMPLE = 16'h3cf3;
		5193: SAMPLE = 16'h3d15;
		5194: SAMPLE = 16'h3d36;
		5195: SAMPLE = 16'h3d57;
		5196: SAMPLE = 16'h3d78;
		5197: SAMPLE = 16'h3d99;
		5198: SAMPLE = 16'h3db9;
		5199: SAMPLE = 16'h3dd8;
		5200: SAMPLE = 16'h3df7;
		5201: SAMPLE = 16'h3e16;
		5202: SAMPLE = 16'h3e34;
		5203: SAMPLE = 16'h3e52;
		5204: SAMPLE = 16'h3e6f;
		5205: SAMPLE = 16'h3e8c;
		5206: SAMPLE = 16'h3ea8;
		5207: SAMPLE = 16'h3ec3;
		5208: SAMPLE = 16'h3ede;
		5209: SAMPLE = 16'h3ef8;
		5210: SAMPLE = 16'h3f11;
		5211: SAMPLE = 16'h3f2a;
		5212: SAMPLE = 16'h3f42;
		5213: SAMPLE = 16'h3f5a;
		5214: SAMPLE = 16'h3f70;
		5215: SAMPLE = 16'h3f86;
		5216: SAMPLE = 16'h3f9b;
		5217: SAMPLE = 16'h3fb0;
		5218: SAMPLE = 16'h3fc4;
		5219: SAMPLE = 16'h3fd6;
		5220: SAMPLE = 16'h3fe8;
		5221: SAMPLE = 16'h3ffa;
		5222: SAMPLE = 16'h400a;
		5223: SAMPLE = 16'h401a;
		5224: SAMPLE = 16'h4029;
		5225: SAMPLE = 16'h4037;
		5226: SAMPLE = 16'h4044;
		5227: SAMPLE = 16'h4050;
		5228: SAMPLE = 16'h405c;
		5229: SAMPLE = 16'h4067;
		5230: SAMPLE = 16'h4071;
		5231: SAMPLE = 16'h407a;
		5232: SAMPLE = 16'h4082;
		5233: SAMPLE = 16'h408a;
		5234: SAMPLE = 16'h4091;
		5235: SAMPLE = 16'h4097;
		5236: SAMPLE = 16'h409c;
		5237: SAMPLE = 16'h40a0;
		5238: SAMPLE = 16'h40a4;
		5239: SAMPLE = 16'h40a7;
		5240: SAMPLE = 16'h40aa;
		5241: SAMPLE = 16'h40ab;
		5242: SAMPLE = 16'h40ac;
		5243: SAMPLE = 16'h40ac;
		5244: SAMPLE = 16'h40ac;
		5245: SAMPLE = 16'h40ab;
		5246: SAMPLE = 16'h40a9;
		5247: SAMPLE = 16'h40a7;
		5248: SAMPLE = 16'h40a4;
		5249: SAMPLE = 16'h40a1;
		5250: SAMPLE = 16'h409d;
		5251: SAMPLE = 16'h4099;
		5252: SAMPLE = 16'h4094;
		5253: SAMPLE = 16'h408f;
		5254: SAMPLE = 16'h4089;
		5255: SAMPLE = 16'h4083;
		5256: SAMPLE = 16'h407c;
		5257: SAMPLE = 16'h4076;
		5258: SAMPLE = 16'h406e;
		5259: SAMPLE = 16'h4067;
		5260: SAMPLE = 16'h405f;
		5261: SAMPLE = 16'h4058;
		5262: SAMPLE = 16'h4050;
		5263: SAMPLE = 16'h4047;
		5264: SAMPLE = 16'h403f;
		5265: SAMPLE = 16'h4037;
		5266: SAMPLE = 16'h402e;
		5267: SAMPLE = 16'h4026;
		5268: SAMPLE = 16'h401d;
		5269: SAMPLE = 16'h4015;
		5270: SAMPLE = 16'h400c;
		5271: SAMPLE = 16'h4004;
		5272: SAMPLE = 16'h3ffc;
		5273: SAMPLE = 16'h3ff4;
		5274: SAMPLE = 16'h3fec;
		5275: SAMPLE = 16'h3fe5;
		5276: SAMPLE = 16'h3fdd;
		5277: SAMPLE = 16'h3fd6;
		5278: SAMPLE = 16'h3fd0;
		5279: SAMPLE = 16'h3fc9;
		5280: SAMPLE = 16'h3fc3;
		5281: SAMPLE = 16'h3fbd;
		5282: SAMPLE = 16'h3fb8;
		5283: SAMPLE = 16'h3fb4;
		5284: SAMPLE = 16'h3faf;
		5285: SAMPLE = 16'h3fac;
		5286: SAMPLE = 16'h3fa8;
		5287: SAMPLE = 16'h3fa6;
		5288: SAMPLE = 16'h3fa4;
		5289: SAMPLE = 16'h3fa2;
		5290: SAMPLE = 16'h3fa2;
		5291: SAMPLE = 16'h3fa2;
		5292: SAMPLE = 16'h3fa2;
		5293: SAMPLE = 16'h3fa3;
		5294: SAMPLE = 16'h3fa5;
		5295: SAMPLE = 16'h3fa8;
		5296: SAMPLE = 16'h3fac;
		5297: SAMPLE = 16'h3fb0;
		5298: SAMPLE = 16'h3fb5;
		5299: SAMPLE = 16'h3fbb;
		5300: SAMPLE = 16'h3fc1;
		5301: SAMPLE = 16'h3fc9;
		5302: SAMPLE = 16'h3fd1;
		5303: SAMPLE = 16'h3fda;
		5304: SAMPLE = 16'h3fe4;
		5305: SAMPLE = 16'h3fef;
		5306: SAMPLE = 16'h3ffb;
		5307: SAMPLE = 16'h4008;
		5308: SAMPLE = 16'h4015;
		5309: SAMPLE = 16'h4024;
		5310: SAMPLE = 16'h4033;
		5311: SAMPLE = 16'h4043;
		5312: SAMPLE = 16'h4054;
		5313: SAMPLE = 16'h4066;
		5314: SAMPLE = 16'h4079;
		5315: SAMPLE = 16'h408d;
		5316: SAMPLE = 16'h40a1;
		5317: SAMPLE = 16'h40b7;
		5318: SAMPLE = 16'h40cd;
		5319: SAMPLE = 16'h40e4;
		5320: SAMPLE = 16'h40fc;
		5321: SAMPLE = 16'h4115;
		5322: SAMPLE = 16'h412e;
		5323: SAMPLE = 16'h4149;
		5324: SAMPLE = 16'h4164;
		5325: SAMPLE = 16'h4180;
		5326: SAMPLE = 16'h419c;
		5327: SAMPLE = 16'h41ba;
		5328: SAMPLE = 16'h41d8;
		5329: SAMPLE = 16'h41f7;
		5330: SAMPLE = 16'h4216;
		5331: SAMPLE = 16'h4236;
		5332: SAMPLE = 16'h4256;
		5333: SAMPLE = 16'h4278;
		5334: SAMPLE = 16'h4299;
		5335: SAMPLE = 16'h42bc;
		5336: SAMPLE = 16'h42de;
		5337: SAMPLE = 16'h4302;
		5338: SAMPLE = 16'h4325;
		5339: SAMPLE = 16'h434a;
		5340: SAMPLE = 16'h436e;
		5341: SAMPLE = 16'h4393;
		5342: SAMPLE = 16'h43b8;
		5343: SAMPLE = 16'h43de;
		5344: SAMPLE = 16'h4403;
		5345: SAMPLE = 16'h4429;
		5346: SAMPLE = 16'h444f;
		5347: SAMPLE = 16'h4476;
		5348: SAMPLE = 16'h449c;
		5349: SAMPLE = 16'h44c3;
		5350: SAMPLE = 16'h44e9;
		5351: SAMPLE = 16'h4510;
		5352: SAMPLE = 16'h4537;
		5353: SAMPLE = 16'h455d;
		5354: SAMPLE = 16'h4584;
		5355: SAMPLE = 16'h45aa;
		5356: SAMPLE = 16'h45d0;
		5357: SAMPLE = 16'h45f6;
		5358: SAMPLE = 16'h461c;
		5359: SAMPLE = 16'h4642;
		5360: SAMPLE = 16'h4667;
		5361: SAMPLE = 16'h468c;
		5362: SAMPLE = 16'h46b0;
		5363: SAMPLE = 16'h46d5;
		5364: SAMPLE = 16'h46f8;
		5365: SAMPLE = 16'h471c;
		5366: SAMPLE = 16'h473f;
		5367: SAMPLE = 16'h4761;
		5368: SAMPLE = 16'h4783;
		5369: SAMPLE = 16'h47a4;
		5370: SAMPLE = 16'h47c5;
		5371: SAMPLE = 16'h47e5;
		5372: SAMPLE = 16'h4804;
		5373: SAMPLE = 16'h4823;
		5374: SAMPLE = 16'h4841;
		5375: SAMPLE = 16'h485e;
		5376: SAMPLE = 16'h487a;
		5377: SAMPLE = 16'h4896;
		5378: SAMPLE = 16'h48b1;
		5379: SAMPLE = 16'h48cb;
		5380: SAMPLE = 16'h48e4;
		5381: SAMPLE = 16'h48fd;
		5382: SAMPLE = 16'h4914;
		5383: SAMPLE = 16'h492b;
		5384: SAMPLE = 16'h4941;
		5385: SAMPLE = 16'h4956;
		5386: SAMPLE = 16'h496a;
		5387: SAMPLE = 16'h497d;
		5388: SAMPLE = 16'h498f;
		5389: SAMPLE = 16'h49a0;
		5390: SAMPLE = 16'h49b0;
		5391: SAMPLE = 16'h49bf;
		5392: SAMPLE = 16'h49cd;
		5393: SAMPLE = 16'h49da;
		5394: SAMPLE = 16'h49e7;
		5395: SAMPLE = 16'h49f2;
		5396: SAMPLE = 16'h49fc;
		5397: SAMPLE = 16'h4a06;
		5398: SAMPLE = 16'h4a0e;
		5399: SAMPLE = 16'h4a16;
		5400: SAMPLE = 16'h4a1c;
		5401: SAMPLE = 16'h4a22;
		5402: SAMPLE = 16'h4a26;
		5403: SAMPLE = 16'h4a2a;
		5404: SAMPLE = 16'h4a2d;
		5405: SAMPLE = 16'h4a2f;
		5406: SAMPLE = 16'h4a30;
		5407: SAMPLE = 16'h4a30;
		5408: SAMPLE = 16'h4a2f;
		5409: SAMPLE = 16'h4a2e;
		5410: SAMPLE = 16'h4a2c;
		5411: SAMPLE = 16'h4a29;
		5412: SAMPLE = 16'h4a25;
		5413: SAMPLE = 16'h4a20;
		5414: SAMPLE = 16'h4a1b;
		5415: SAMPLE = 16'h4a15;
		5416: SAMPLE = 16'h4a0e;
		5417: SAMPLE = 16'h4a07;
		5418: SAMPLE = 16'h49ff;
		5419: SAMPLE = 16'h49f7;
		5420: SAMPLE = 16'h49ee;
		5421: SAMPLE = 16'h49e4;
		5422: SAMPLE = 16'h49da;
		5423: SAMPLE = 16'h49d0;
		5424: SAMPLE = 16'h49c5;
		5425: SAMPLE = 16'h49ba;
		5426: SAMPLE = 16'h49ae;
		5427: SAMPLE = 16'h49a2;
		5428: SAMPLE = 16'h4996;
		5429: SAMPLE = 16'h498a;
		5430: SAMPLE = 16'h497d;
		5431: SAMPLE = 16'h4970;
		5432: SAMPLE = 16'h4963;
		5433: SAMPLE = 16'h4956;
		5434: SAMPLE = 16'h4949;
		5435: SAMPLE = 16'h493c;
		5436: SAMPLE = 16'h492f;
		5437: SAMPLE = 16'h4922;
		5438: SAMPLE = 16'h4915;
		5439: SAMPLE = 16'h4909;
		5440: SAMPLE = 16'h48fc;
		5441: SAMPLE = 16'h48f0;
		5442: SAMPLE = 16'h48e4;
		5443: SAMPLE = 16'h48d8;
		5444: SAMPLE = 16'h48cc;
		5445: SAMPLE = 16'h48c1;
		5446: SAMPLE = 16'h48b6;
		5447: SAMPLE = 16'h48ac;
		5448: SAMPLE = 16'h48a2;
		5449: SAMPLE = 16'h4899;
		5450: SAMPLE = 16'h4890;
		5451: SAMPLE = 16'h4888;
		5452: SAMPLE = 16'h4881;
		5453: SAMPLE = 16'h487a;
		5454: SAMPLE = 16'h4873;
		5455: SAMPLE = 16'h486e;
		5456: SAMPLE = 16'h4869;
		5457: SAMPLE = 16'h4865;
		5458: SAMPLE = 16'h4862;
		5459: SAMPLE = 16'h485f;
		5460: SAMPLE = 16'h485e;
		5461: SAMPLE = 16'h485d;
		5462: SAMPLE = 16'h485d;
		5463: SAMPLE = 16'h485e;
		5464: SAMPLE = 16'h4860;
		5465: SAMPLE = 16'h4863;
		5466: SAMPLE = 16'h4867;
		5467: SAMPLE = 16'h486c;
		5468: SAMPLE = 16'h4872;
		5469: SAMPLE = 16'h4879;
		5470: SAMPLE = 16'h4881;
		5471: SAMPLE = 16'h488a;
		5472: SAMPLE = 16'h4894;
		5473: SAMPLE = 16'h489f;
		5474: SAMPLE = 16'h48ab;
		5475: SAMPLE = 16'h48b8;
		5476: SAMPLE = 16'h48c7;
		5477: SAMPLE = 16'h48d6;
		5478: SAMPLE = 16'h48e6;
		5479: SAMPLE = 16'h48f8;
		5480: SAMPLE = 16'h490b;
		5481: SAMPLE = 16'h491e;
		5482: SAMPLE = 16'h4933;
		5483: SAMPLE = 16'h4949;
		5484: SAMPLE = 16'h4960;
		5485: SAMPLE = 16'h4978;
		5486: SAMPLE = 16'h4990;
		5487: SAMPLE = 16'h49aa;
		5488: SAMPLE = 16'h49c5;
		5489: SAMPLE = 16'h49e1;
		5490: SAMPLE = 16'h49fe;
		5491: SAMPLE = 16'h4a1c;
		5492: SAMPLE = 16'h4a3b;
		5493: SAMPLE = 16'h4a5b;
		5494: SAMPLE = 16'h4a7b;
		5495: SAMPLE = 16'h4a9d;
		5496: SAMPLE = 16'h4abf;
		5497: SAMPLE = 16'h4ae2;
		5498: SAMPLE = 16'h4b06;
		5499: SAMPLE = 16'h4b2b;
		5500: SAMPLE = 16'h4b51;
		5501: SAMPLE = 16'h4b77;
		5502: SAMPLE = 16'h4b9e;
		5503: SAMPLE = 16'h4bc5;
		5504: SAMPLE = 16'h4bed;
		5505: SAMPLE = 16'h4c16;
		5506: SAMPLE = 16'h4c3f;
		5507: SAMPLE = 16'h4c68;
		5508: SAMPLE = 16'h4c93;
		5509: SAMPLE = 16'h4cbd;
		5510: SAMPLE = 16'h4ce8;
		5511: SAMPLE = 16'h4d13;
		5512: SAMPLE = 16'h4d3f;
		5513: SAMPLE = 16'h4d6a;
		5514: SAMPLE = 16'h4d96;
		5515: SAMPLE = 16'h4dc3;
		5516: SAMPLE = 16'h4def;
		5517: SAMPLE = 16'h4e1b;
		5518: SAMPLE = 16'h4e48;
		5519: SAMPLE = 16'h4e74;
		5520: SAMPLE = 16'h4ea1;
		5521: SAMPLE = 16'h4ecd;
		5522: SAMPLE = 16'h4ef9;
		5523: SAMPLE = 16'h4f25;
		5524: SAMPLE = 16'h4f51;
		5525: SAMPLE = 16'h4f7d;
		5526: SAMPLE = 16'h4fa8;
		5527: SAMPLE = 16'h4fd3;
		5528: SAMPLE = 16'h4ffd;
		5529: SAMPLE = 16'h5027;
		5530: SAMPLE = 16'h5051;
		5531: SAMPLE = 16'h507a;
		5532: SAMPLE = 16'h50a3;
		5533: SAMPLE = 16'h50cb;
		5534: SAMPLE = 16'h50f2;
		5535: SAMPLE = 16'h5119;
		5536: SAMPLE = 16'h513f;
		5537: SAMPLE = 16'h5165;
		5538: SAMPLE = 16'h5189;
		5539: SAMPLE = 16'h51ad;
		5540: SAMPLE = 16'h51d0;
		5541: SAMPLE = 16'h51f2;
		5542: SAMPLE = 16'h5213;
		5543: SAMPLE = 16'h5233;
		5544: SAMPLE = 16'h5253;
		5545: SAMPLE = 16'h5271;
		5546: SAMPLE = 16'h528e;
		5547: SAMPLE = 16'h52ab;
		5548: SAMPLE = 16'h52c6;
		5549: SAMPLE = 16'h52e0;
		5550: SAMPLE = 16'h52f9;
		5551: SAMPLE = 16'h5311;
		5552: SAMPLE = 16'h5328;
		5553: SAMPLE = 16'h533d;
		5554: SAMPLE = 16'h5352;
		5555: SAMPLE = 16'h5365;
		5556: SAMPLE = 16'h5377;
		5557: SAMPLE = 16'h5388;
		5558: SAMPLE = 16'h5398;
		5559: SAMPLE = 16'h53a6;
		5560: SAMPLE = 16'h53b4;
		5561: SAMPLE = 16'h53c0;
		5562: SAMPLE = 16'h53ca;
		5563: SAMPLE = 16'h53d4;
		5564: SAMPLE = 16'h53dc;
		5565: SAMPLE = 16'h53e4;
		5566: SAMPLE = 16'h53ea;
		5567: SAMPLE = 16'h53ee;
		5568: SAMPLE = 16'h53f2;
		5569: SAMPLE = 16'h53f4;
		5570: SAMPLE = 16'h53f6;
		5571: SAMPLE = 16'h53f6;
		5572: SAMPLE = 16'h53f5;
		5573: SAMPLE = 16'h53f2;
		5574: SAMPLE = 16'h53ef;
		5575: SAMPLE = 16'h53eb;
		5576: SAMPLE = 16'h53e5;
		5577: SAMPLE = 16'h53df;
		5578: SAMPLE = 16'h53d7;
		5579: SAMPLE = 16'h53cf;
		5580: SAMPLE = 16'h53c6;
		5581: SAMPLE = 16'h53bb;
		5582: SAMPLE = 16'h53b0;
		5583: SAMPLE = 16'h53a4;
		5584: SAMPLE = 16'h5397;
		5585: SAMPLE = 16'h5389;
		5586: SAMPLE = 16'h537b;
		5587: SAMPLE = 16'h536c;
		5588: SAMPLE = 16'h535c;
		5589: SAMPLE = 16'h534b;
		5590: SAMPLE = 16'h533a;
		5591: SAMPLE = 16'h5329;
		5592: SAMPLE = 16'h5317;
		5593: SAMPLE = 16'h5304;
		5594: SAMPLE = 16'h52f1;
		5595: SAMPLE = 16'h52de;
		5596: SAMPLE = 16'h52ca;
		5597: SAMPLE = 16'h52b6;
		5598: SAMPLE = 16'h52a2;
		5599: SAMPLE = 16'h528d;
		5600: SAMPLE = 16'h5279;
		5601: SAMPLE = 16'h5264;
		5602: SAMPLE = 16'h524f;
		5603: SAMPLE = 16'h523b;
		5604: SAMPLE = 16'h5226;
		5605: SAMPLE = 16'h5212;
		5606: SAMPLE = 16'h51fd;
		5607: SAMPLE = 16'h51e9;
		5608: SAMPLE = 16'h51d5;
		5609: SAMPLE = 16'h51c2;
		5610: SAMPLE = 16'h51ae;
		5611: SAMPLE = 16'h519b;
		5612: SAMPLE = 16'h5189;
		5613: SAMPLE = 16'h5177;
		5614: SAMPLE = 16'h5166;
		5615: SAMPLE = 16'h5155;
		5616: SAMPLE = 16'h5145;
		5617: SAMPLE = 16'h5135;
		5618: SAMPLE = 16'h5126;
		5619: SAMPLE = 16'h5118;
		5620: SAMPLE = 16'h510b;
		5621: SAMPLE = 16'h50ff;
		5622: SAMPLE = 16'h50f3;
		5623: SAMPLE = 16'h50e9;
		5624: SAMPLE = 16'h50df;
		5625: SAMPLE = 16'h50d7;
		5626: SAMPLE = 16'h50cf;
		5627: SAMPLE = 16'h50c9;
		5628: SAMPLE = 16'h50c3;
		5629: SAMPLE = 16'h50bf;
		5630: SAMPLE = 16'h50bc;
		5631: SAMPLE = 16'h50ba;
		5632: SAMPLE = 16'h50ba;
		5633: SAMPLE = 16'h50ba;
		5634: SAMPLE = 16'h50bc;
		5635: SAMPLE = 16'h50bf;
		5636: SAMPLE = 16'h50c4;
		5637: SAMPLE = 16'h50ca;
		5638: SAMPLE = 16'h50d1;
		5639: SAMPLE = 16'h50d9;
		5640: SAMPLE = 16'h50e3;
		5641: SAMPLE = 16'h50ef;
		5642: SAMPLE = 16'h50fb;
		5643: SAMPLE = 16'h510a;
		5644: SAMPLE = 16'h5119;
		5645: SAMPLE = 16'h512a;
		5646: SAMPLE = 16'h513c;
		5647: SAMPLE = 16'h5150;
		5648: SAMPLE = 16'h5165;
		5649: SAMPLE = 16'h517c;
		5650: SAMPLE = 16'h5194;
		5651: SAMPLE = 16'h51ad;
		5652: SAMPLE = 16'h51c8;
		5653: SAMPLE = 16'h51e4;
		5654: SAMPLE = 16'h5202;
		5655: SAMPLE = 16'h5221;
		5656: SAMPLE = 16'h5241;
		5657: SAMPLE = 16'h5262;
		5658: SAMPLE = 16'h5285;
		5659: SAMPLE = 16'h52a9;
		5660: SAMPLE = 16'h52ce;
		5661: SAMPLE = 16'h52f4;
		5662: SAMPLE = 16'h531c;
		5663: SAMPLE = 16'h5345;
		5664: SAMPLE = 16'h536e;
		5665: SAMPLE = 16'h5399;
		5666: SAMPLE = 16'h53c5;
		5667: SAMPLE = 16'h53f2;
		5668: SAMPLE = 16'h5420;
		5669: SAMPLE = 16'h544f;
		5670: SAMPLE = 16'h547e;
		5671: SAMPLE = 16'h54af;
		5672: SAMPLE = 16'h54e0;
		5673: SAMPLE = 16'h5512;
		5674: SAMPLE = 16'h5544;
		5675: SAMPLE = 16'h5578;
		5676: SAMPLE = 16'h55ac;
		5677: SAMPLE = 16'h55e0;
		5678: SAMPLE = 16'h5615;
		5679: SAMPLE = 16'h564a;
		5680: SAMPLE = 16'h5680;
		5681: SAMPLE = 16'h56b6;
		5682: SAMPLE = 16'h56ec;
		5683: SAMPLE = 16'h5723;
		5684: SAMPLE = 16'h5759;
		5685: SAMPLE = 16'h5790;
		5686: SAMPLE = 16'h57c7;
		5687: SAMPLE = 16'h57fe;
		5688: SAMPLE = 16'h5834;
		5689: SAMPLE = 16'h586b;
		5690: SAMPLE = 16'h58a1;
		5691: SAMPLE = 16'h58d7;
		5692: SAMPLE = 16'h590d;
		5693: SAMPLE = 16'h5943;
		5694: SAMPLE = 16'h5978;
		5695: SAMPLE = 16'h59ac;
		5696: SAMPLE = 16'h59e0;
		5697: SAMPLE = 16'h5a14;
		5698: SAMPLE = 16'h5a47;
		5699: SAMPLE = 16'h5a79;
		5700: SAMPLE = 16'h5aaa;
		5701: SAMPLE = 16'h5adb;
		5702: SAMPLE = 16'h5b0a;
		5703: SAMPLE = 16'h5b39;
		5704: SAMPLE = 16'h5b67;
		5705: SAMPLE = 16'h5b94;
		5706: SAMPLE = 16'h5bc0;
		5707: SAMPLE = 16'h5bea;
		5708: SAMPLE = 16'h5c14;
		5709: SAMPLE = 16'h5c3c;
		5710: SAMPLE = 16'h5c63;
		5711: SAMPLE = 16'h5c89;
		5712: SAMPLE = 16'h5cad;
		5713: SAMPLE = 16'h5cd0;
		5714: SAMPLE = 16'h5cf2;
		5715: SAMPLE = 16'h5d12;
		5716: SAMPLE = 16'h5d31;
		5717: SAMPLE = 16'h5d4f;
		5718: SAMPLE = 16'h5d6a;
		5719: SAMPLE = 16'h5d85;
		5720: SAMPLE = 16'h5d9e;
		5721: SAMPLE = 16'h5db5;
		5722: SAMPLE = 16'h5dca;
		5723: SAMPLE = 16'h5dde;
		5724: SAMPLE = 16'h5df0;
		5725: SAMPLE = 16'h5e01;
		5726: SAMPLE = 16'h5e10;
		5727: SAMPLE = 16'h5e1d;
		5728: SAMPLE = 16'h5e29;
		5729: SAMPLE = 16'h5e33;
		5730: SAMPLE = 16'h5e3b;
		5731: SAMPLE = 16'h5e42;
		5732: SAMPLE = 16'h5e46;
		5733: SAMPLE = 16'h5e4a;
		5734: SAMPLE = 16'h5e4b;
		5735: SAMPLE = 16'h5e4b;
		5736: SAMPLE = 16'h5e49;
		5737: SAMPLE = 16'h5e46;
		5738: SAMPLE = 16'h5e41;
		5739: SAMPLE = 16'h5e3a;
		5740: SAMPLE = 16'h5e32;
		5741: SAMPLE = 16'h5e28;
		5742: SAMPLE = 16'h5e1d;
		5743: SAMPLE = 16'h5e10;
		5744: SAMPLE = 16'h5e01;
		5745: SAMPLE = 16'h5df2;
		5746: SAMPLE = 16'h5de1;
		5747: SAMPLE = 16'h5dce;
		5748: SAMPLE = 16'h5dba;
		5749: SAMPLE = 16'h5da5;
		5750: SAMPLE = 16'h5d8f;
		5751: SAMPLE = 16'h5d77;
		5752: SAMPLE = 16'h5d5f;
		5753: SAMPLE = 16'h5d45;
		5754: SAMPLE = 16'h5d2a;
		5755: SAMPLE = 16'h5d0e;
		5756: SAMPLE = 16'h5cf1;
		5757: SAMPLE = 16'h5cd4;
		5758: SAMPLE = 16'h5cb5;
		5759: SAMPLE = 16'h5c96;
		5760: SAMPLE = 16'h5c76;
		5761: SAMPLE = 16'h5c56;
		5762: SAMPLE = 16'h5c34;
		5763: SAMPLE = 16'h5c13;
		5764: SAMPLE = 16'h5bf1;
		5765: SAMPLE = 16'h5bce;
		5766: SAMPLE = 16'h5bab;
		5767: SAMPLE = 16'h5b88;
		5768: SAMPLE = 16'h5b65;
		5769: SAMPLE = 16'h5b41;
		5770: SAMPLE = 16'h5b1e;
		5771: SAMPLE = 16'h5afb;
		5772: SAMPLE = 16'h5ad7;
		5773: SAMPLE = 16'h5ab4;
		5774: SAMPLE = 16'h5a91;
		5775: SAMPLE = 16'h5a6e;
		5776: SAMPLE = 16'h5a4c;
		5777: SAMPLE = 16'h5a2a;
		5778: SAMPLE = 16'h5a09;
		5779: SAMPLE = 16'h59e8;
		5780: SAMPLE = 16'h59c8;
		5781: SAMPLE = 16'h59a9;
		5782: SAMPLE = 16'h598b;
		5783: SAMPLE = 16'h596d;
		5784: SAMPLE = 16'h5950;
		5785: SAMPLE = 16'h5934;
		5786: SAMPLE = 16'h591a;
		5787: SAMPLE = 16'h5900;
		5788: SAMPLE = 16'h58e8;
		5789: SAMPLE = 16'h58d0;
		5790: SAMPLE = 16'h58bb;
		5791: SAMPLE = 16'h58a6;
		5792: SAMPLE = 16'h5893;
		5793: SAMPLE = 16'h5881;
		5794: SAMPLE = 16'h5871;
		5795: SAMPLE = 16'h5863;
		5796: SAMPLE = 16'h5856;
		5797: SAMPLE = 16'h584b;
		5798: SAMPLE = 16'h5841;
		5799: SAMPLE = 16'h5839;
		5800: SAMPLE = 16'h5833;
		5801: SAMPLE = 16'h582f;
		5802: SAMPLE = 16'h582d;
		5803: SAMPLE = 16'h582d;
		5804: SAMPLE = 16'h582e;
		5805: SAMPLE = 16'h5832;
		5806: SAMPLE = 16'h5838;
		5807: SAMPLE = 16'h583f;
		5808: SAMPLE = 16'h5849;
		5809: SAMPLE = 16'h5855;
		5810: SAMPLE = 16'h5862;
		5811: SAMPLE = 16'h5872;
		5812: SAMPLE = 16'h5884;
		5813: SAMPLE = 16'h5898;
		5814: SAMPLE = 16'h58ae;
		5815: SAMPLE = 16'h58c7;
		5816: SAMPLE = 16'h58e1;
		5817: SAMPLE = 16'h58fe;
		5818: SAMPLE = 16'h591c;
		5819: SAMPLE = 16'h593d;
		5820: SAMPLE = 16'h595f;
		5821: SAMPLE = 16'h5984;
		5822: SAMPLE = 16'h59ab;
		5823: SAMPLE = 16'h59d4;
		5824: SAMPLE = 16'h59ff;
		5825: SAMPLE = 16'h5a2b;
		5826: SAMPLE = 16'h5a5a;
		5827: SAMPLE = 16'h5a8b;
		5828: SAMPLE = 16'h5abd;
		5829: SAMPLE = 16'h5af1;
		5830: SAMPLE = 16'h5b27;
		5831: SAMPLE = 16'h5b5f;
		5832: SAMPLE = 16'h5b98;
		5833: SAMPLE = 16'h5bd3;
		5834: SAMPLE = 16'h5c10;
		5835: SAMPLE = 16'h5c4e;
		5836: SAMPLE = 16'h5c8e;
		5837: SAMPLE = 16'h5ccf;
		5838: SAMPLE = 16'h5d11;
		5839: SAMPLE = 16'h5d55;
		5840: SAMPLE = 16'h5d99;
		5841: SAMPLE = 16'h5ddf;
		5842: SAMPLE = 16'h5e26;
		5843: SAMPLE = 16'h5e6e;
		5844: SAMPLE = 16'h5eb7;
		5845: SAMPLE = 16'h5f01;
		5846: SAMPLE = 16'h5f4b;
		5847: SAMPLE = 16'h5f96;
		5848: SAMPLE = 16'h5fe2;
		5849: SAMPLE = 16'h602e;
		5850: SAMPLE = 16'h607b;
		5851: SAMPLE = 16'h60c8;
		5852: SAMPLE = 16'h6115;
		5853: SAMPLE = 16'h6162;
		5854: SAMPLE = 16'h61b0;
		5855: SAMPLE = 16'h61fd;
		5856: SAMPLE = 16'h624a;
		5857: SAMPLE = 16'h6297;
		5858: SAMPLE = 16'h62e4;
		5859: SAMPLE = 16'h6331;
		5860: SAMPLE = 16'h637d;
		5861: SAMPLE = 16'h63c8;
		5862: SAMPLE = 16'h6413;
		5863: SAMPLE = 16'h645d;
		5864: SAMPLE = 16'h64a6;
		5865: SAMPLE = 16'h64ee;
		5866: SAMPLE = 16'h6536;
		5867: SAMPLE = 16'h657c;
		5868: SAMPLE = 16'h65c1;
		5869: SAMPLE = 16'h6605;
		5870: SAMPLE = 16'h6647;
		5871: SAMPLE = 16'h6688;
		5872: SAMPLE = 16'h66c7;
		5873: SAMPLE = 16'h6705;
		5874: SAMPLE = 16'h6741;
		5875: SAMPLE = 16'h677c;
		5876: SAMPLE = 16'h67b4;
		5877: SAMPLE = 16'h67eb;
		5878: SAMPLE = 16'h681f;
		5879: SAMPLE = 16'h6852;
		5880: SAMPLE = 16'h6882;
		5881: SAMPLE = 16'h68b1;
		5882: SAMPLE = 16'h68dd;
		5883: SAMPLE = 16'h6906;
		5884: SAMPLE = 16'h692e;
		5885: SAMPLE = 16'h6953;
		5886: SAMPLE = 16'h6975;
		5887: SAMPLE = 16'h6995;
		5888: SAMPLE = 16'h69b2;
		5889: SAMPLE = 16'h69cd;
		5890: SAMPLE = 16'h69e5;
		5891: SAMPLE = 16'h69fb;
		5892: SAMPLE = 16'h6a0e;
		5893: SAMPLE = 16'h6a1e;
		5894: SAMPLE = 16'h6a2b;
		5895: SAMPLE = 16'h6a35;
		5896: SAMPLE = 16'h6a3d;
		5897: SAMPLE = 16'h6a42;
		5898: SAMPLE = 16'h6a44;
		5899: SAMPLE = 16'h6a43;
		5900: SAMPLE = 16'h6a40;
		5901: SAMPLE = 16'h6a39;
		5902: SAMPLE = 16'h6a30;
		5903: SAMPLE = 16'h6a24;
		5904: SAMPLE = 16'h6a15;
		5905: SAMPLE = 16'h6a04;
		5906: SAMPLE = 16'h69f0;
		5907: SAMPLE = 16'h69d8;
		5908: SAMPLE = 16'h69bf;
		5909: SAMPLE = 16'h69a2;
		5910: SAMPLE = 16'h6983;
		5911: SAMPLE = 16'h6962;
		5912: SAMPLE = 16'h693d;
		5913: SAMPLE = 16'h6917;
		5914: SAMPLE = 16'h68ee;
		5915: SAMPLE = 16'h68c2;
		5916: SAMPLE = 16'h6894;
		5917: SAMPLE = 16'h6864;
		5918: SAMPLE = 16'h6832;
		5919: SAMPLE = 16'h67fe;
		5920: SAMPLE = 16'h67c7;
		5921: SAMPLE = 16'h678f;
		5922: SAMPLE = 16'h6755;
		5923: SAMPLE = 16'h6719;
		5924: SAMPLE = 16'h66db;
		5925: SAMPLE = 16'h669c;
		5926: SAMPLE = 16'h665b;
		5927: SAMPLE = 16'h6619;
		5928: SAMPLE = 16'h65d5;
		5929: SAMPLE = 16'h6590;
		5930: SAMPLE = 16'h654a;
		5931: SAMPLE = 16'h6503;
		5932: SAMPLE = 16'h64bc;
		5933: SAMPLE = 16'h6473;
		5934: SAMPLE = 16'h642a;
		5935: SAMPLE = 16'h63e0;
		5936: SAMPLE = 16'h6396;
		5937: SAMPLE = 16'h634c;
		5938: SAMPLE = 16'h6301;
		5939: SAMPLE = 16'h62b6;
		5940: SAMPLE = 16'h626c;
		5941: SAMPLE = 16'h6221;
		5942: SAMPLE = 16'h61d7;
		5943: SAMPLE = 16'h618d;
		5944: SAMPLE = 16'h6144;
		5945: SAMPLE = 16'h60fc;
		5946: SAMPLE = 16'h60b4;
		5947: SAMPLE = 16'h606e;
		5948: SAMPLE = 16'h6029;
		5949: SAMPLE = 16'h5fe4;
		5950: SAMPLE = 16'h5fa2;
		5951: SAMPLE = 16'h5f60;
		5952: SAMPLE = 16'h5f20;
		5953: SAMPLE = 16'h5ee3;
		5954: SAMPLE = 16'h5ea6;
		5955: SAMPLE = 16'h5e6c;
		5956: SAMPLE = 16'h5e34;
		5957: SAMPLE = 16'h5dff;
		5958: SAMPLE = 16'h5dcb;
		5959: SAMPLE = 16'h5d9a;
		5960: SAMPLE = 16'h5d6c;
		5961: SAMPLE = 16'h5d40;
		5962: SAMPLE = 16'h5d18;
		5963: SAMPLE = 16'h5cf2;
		5964: SAMPLE = 16'h5ccf;
		5965: SAMPLE = 16'h5caf;
		5966: SAMPLE = 16'h5c93;
		5967: SAMPLE = 16'h5c7a;
		5968: SAMPLE = 16'h5c64;
		5969: SAMPLE = 16'h5c52;
		5970: SAMPLE = 16'h5c44;
		5971: SAMPLE = 16'h5c39;
		5972: SAMPLE = 16'h5c32;
		5973: SAMPLE = 16'h5c2e;
		5974: SAMPLE = 16'h5c2f;
		5975: SAMPLE = 16'h5c34;
		5976: SAMPLE = 16'h5c3c;
		5977: SAMPLE = 16'h5c49;
		5978: SAMPLE = 16'h5c5a;
		5979: SAMPLE = 16'h5c6f;
		5980: SAMPLE = 16'h5c88;
		5981: SAMPLE = 16'h5ca6;
		5982: SAMPLE = 16'h5cc8;
		5983: SAMPLE = 16'h5cee;
		5984: SAMPLE = 16'h5d18;
		5985: SAMPLE = 16'h5d47;
		5986: SAMPLE = 16'h5d7a;
		5987: SAMPLE = 16'h5db2;
		5988: SAMPLE = 16'h5dee;
		5989: SAMPLE = 16'h5e2e;
		5990: SAMPLE = 16'h5e73;
		5991: SAMPLE = 16'h5ebc;
		5992: SAMPLE = 16'h5f09;
		5993: SAMPLE = 16'h5f5a;
		5994: SAMPLE = 16'h5fb0;
		5995: SAMPLE = 16'h600a;
		5996: SAMPLE = 16'h6067;
		5997: SAMPLE = 16'h60c9;
		5998: SAMPLE = 16'h612f;
		5999: SAMPLE = 16'h6199;
		6000: SAMPLE = 16'h6207;
		6001: SAMPLE = 16'h6278;
		6002: SAMPLE = 16'h62ee;
		6003: SAMPLE = 16'h6366;
		6004: SAMPLE = 16'h63e2;
		6005: SAMPLE = 16'h6462;
		6006: SAMPLE = 16'h64e5;
		6007: SAMPLE = 16'h656b;
		6008: SAMPLE = 16'h65f4;
		6009: SAMPLE = 16'h667f;
		6010: SAMPLE = 16'h670e;
		6011: SAMPLE = 16'h679f;
		6012: SAMPLE = 16'h6833;
		6013: SAMPLE = 16'h68c9;
		6014: SAMPLE = 16'h6961;
		6015: SAMPLE = 16'h69fb;
		6016: SAMPLE = 16'h6a97;
		6017: SAMPLE = 16'h6b34;
		6018: SAMPLE = 16'h6bd3;
		6019: SAMPLE = 16'h6c73;
		6020: SAMPLE = 16'h6d15;
		6021: SAMPLE = 16'h6db7;
		6022: SAMPLE = 16'h6e5a;
		6023: SAMPLE = 16'h6efd;
		6024: SAMPLE = 16'h6fa1;
		6025: SAMPLE = 16'h7045;
		6026: SAMPLE = 16'h70e9;
		6027: SAMPLE = 16'h718c;
		6028: SAMPLE = 16'h722f;
		6029: SAMPLE = 16'h72d1;
		6030: SAMPLE = 16'h7372;
		6031: SAMPLE = 16'h7412;
		6032: SAMPLE = 16'h74b0;
		6033: SAMPLE = 16'h754d;
		6034: SAMPLE = 16'h75e7;
		6035: SAMPLE = 16'h7680;
		6036: SAMPLE = 16'h7716;
		6037: SAMPLE = 16'h77aa;
		6038: SAMPLE = 16'h783a;
		6039: SAMPLE = 16'h78c8;
		6040: SAMPLE = 16'h7952;
		6041: SAMPLE = 16'h79d8;
		6042: SAMPLE = 16'h7a5b;
		6043: SAMPLE = 16'h7ada;
		6044: SAMPLE = 16'h7b54;
		6045: SAMPLE = 16'h7bca;
		6046: SAMPLE = 16'h7c3b;
		6047: SAMPLE = 16'h7ca7;
		6048: SAMPLE = 16'h7d0e;
		6049: SAMPLE = 16'h7d6f;
		6050: SAMPLE = 16'h7dca;
		6051: SAMPLE = 16'h7e1f;
		6052: SAMPLE = 16'h7e6f;
		6053: SAMPLE = 16'h7eb7;
		6054: SAMPLE = 16'h7ef9;
		6055: SAMPLE = 16'h7f35;
		6056: SAMPLE = 16'h7f69;
		6057: SAMPLE = 16'h7f95;
		6058: SAMPLE = 16'h7fba;
		6059: SAMPLE = 16'h7fd8;
		6060: SAMPLE = 16'h7fed;
		6061: SAMPLE = 16'h7ffb;
		6062: SAMPLE = 16'h8000;
		6063: SAMPLE = 16'h7ffc;
		6064: SAMPLE = 16'h7ff0;
		6065: SAMPLE = 16'h7fda;
		6066: SAMPLE = 16'h7fbc;
		6067: SAMPLE = 16'h7f94;
		6068: SAMPLE = 16'h7f63;
		6069: SAMPLE = 16'h7f29;
		6070: SAMPLE = 16'h7ee4;
		6071: SAMPLE = 16'h7e96;
		6072: SAMPLE = 16'h7e3e;
		6073: SAMPLE = 16'h7ddb;
		6074: SAMPLE = 16'h7d6e;
		6075: SAMPLE = 16'h7cf7;
		6076: SAMPLE = 16'h7c75;
		6077: SAMPLE = 16'h7be9;
		6078: SAMPLE = 16'h7b52;
		6079: SAMPLE = 16'h7ab0;
		6080: SAMPLE = 16'h7a03;
		6081: SAMPLE = 16'h794c;
		6082: SAMPLE = 16'h7889;
		6083: SAMPLE = 16'h77bb;
		6084: SAMPLE = 16'h76e2;
		6085: SAMPLE = 16'h75fe;
		6086: SAMPLE = 16'h750e;
		6087: SAMPLE = 16'h7413;
		6088: SAMPLE = 16'h730d;
		6089: SAMPLE = 16'h71fc;
		6090: SAMPLE = 16'h70df;
		6091: SAMPLE = 16'h6fb8;
		6092: SAMPLE = 16'h6e84;
		6093: SAMPLE = 16'h6d46;
		6094: SAMPLE = 16'h6bfd;
		6095: SAMPLE = 16'h6aa8;
		6096: SAMPLE = 16'h6948;
		6097: SAMPLE = 16'h67dd;
		6098: SAMPLE = 16'h6667;
		6099: SAMPLE = 16'h64e6;
		6100: SAMPLE = 16'h635b;
		6101: SAMPLE = 16'h61c5;
		6102: SAMPLE = 16'h6024;
		6103: SAMPLE = 16'h5e78;
		6104: SAMPLE = 16'h5cc2;
		6105: SAMPLE = 16'h5b02;
		6106: SAMPLE = 16'h5938;
		6107: SAMPLE = 16'h5764;
		6108: SAMPLE = 16'h5586;
		6109: SAMPLE = 16'h539e;
		6110: SAMPLE = 16'h51ad;
		6111: SAMPLE = 16'h4fb3;
		6112: SAMPLE = 16'h4daf;
		6113: SAMPLE = 16'h4ba2;
		6114: SAMPLE = 16'h498d;
		6115: SAMPLE = 16'h476f;
		6116: SAMPLE = 16'h4549;
		6117: SAMPLE = 16'h431b;
		6118: SAMPLE = 16'h40e5;
		6119: SAMPLE = 16'h3ea7;
		6120: SAMPLE = 16'h3c62;
		6121: SAMPLE = 16'h3a15;
		6122: SAMPLE = 16'h37c2;
		6123: SAMPLE = 16'h3568;
		6124: SAMPLE = 16'h3308;
		6125: SAMPLE = 16'h30a1;
		6126: SAMPLE = 16'h2e35;
		6127: SAMPLE = 16'h2bc3;
		6128: SAMPLE = 16'h294c;
		6129: SAMPLE = 16'h26d0;
		6130: SAMPLE = 16'h244f;
		6131: SAMPLE = 16'h21ca;
		6132: SAMPLE = 16'h1f40;
		6133: SAMPLE = 16'h1cb3;
		6134: SAMPLE = 16'h1a22;
		6135: SAMPLE = 16'h178e;
		6136: SAMPLE = 16'h14f7;
		6137: SAMPLE = 16'h125e;
		6138: SAMPLE = 16'hfc3;
		6139: SAMPLE = 16'hd25;
		6140: SAMPLE = 16'ha86;
		6141: SAMPLE = 16'h7e5;
		6142: SAMPLE = 16'h544;
		6143: SAMPLE = 16'h2a2;
		6144: SAMPLE = 16'h0;
		6145: SAMPLE = 16'hfd5d;
		6146: SAMPLE = 16'hfabb;
		6147: SAMPLE = 16'hf81a;
		6148: SAMPLE = 16'hf579;
		6149: SAMPLE = 16'hf2da;
		6150: SAMPLE = 16'hf03c;
		6151: SAMPLE = 16'heda1;
		6152: SAMPLE = 16'heb08;
		6153: SAMPLE = 16'he871;
		6154: SAMPLE = 16'he5dd;
		6155: SAMPLE = 16'he34c;
		6156: SAMPLE = 16'he0bf;
		6157: SAMPLE = 16'hde35;
		6158: SAMPLE = 16'hdbb0;
		6159: SAMPLE = 16'hd92f;
		6160: SAMPLE = 16'hd6b3;
		6161: SAMPLE = 16'hd43c;
		6162: SAMPLE = 16'hd1ca;
		6163: SAMPLE = 16'hcf5e;
		6164: SAMPLE = 16'hccf7;
		6165: SAMPLE = 16'hca97;
		6166: SAMPLE = 16'hc83d;
		6167: SAMPLE = 16'hc5ea;
		6168: SAMPLE = 16'hc39d;
		6169: SAMPLE = 16'hc158;
		6170: SAMPLE = 16'hbf1a;
		6171: SAMPLE = 16'hbce4;
		6172: SAMPLE = 16'hbab6;
		6173: SAMPLE = 16'hb890;
		6174: SAMPLE = 16'hb672;
		6175: SAMPLE = 16'hb45d;
		6176: SAMPLE = 16'hb250;
		6177: SAMPLE = 16'hb04c;
		6178: SAMPLE = 16'hae52;
		6179: SAMPLE = 16'hac61;
		6180: SAMPLE = 16'haa79;
		6181: SAMPLE = 16'ha89b;
		6182: SAMPLE = 16'ha6c7;
		6183: SAMPLE = 16'ha4fd;
		6184: SAMPLE = 16'ha33d;
		6185: SAMPLE = 16'ha187;
		6186: SAMPLE = 16'h9fdb;
		6187: SAMPLE = 16'h9e3a;
		6188: SAMPLE = 16'h9ca4;
		6189: SAMPLE = 16'h9b19;
		6190: SAMPLE = 16'h9998;
		6191: SAMPLE = 16'h9822;
		6192: SAMPLE = 16'h96b7;
		6193: SAMPLE = 16'h9557;
		6194: SAMPLE = 16'h9402;
		6195: SAMPLE = 16'h92b9;
		6196: SAMPLE = 16'h917b;
		6197: SAMPLE = 16'h9047;
		6198: SAMPLE = 16'h8f20;
		6199: SAMPLE = 16'h8e03;
		6200: SAMPLE = 16'h8cf2;
		6201: SAMPLE = 16'h8bec;
		6202: SAMPLE = 16'h8af1;
		6203: SAMPLE = 16'h8a01;
		6204: SAMPLE = 16'h891d;
		6205: SAMPLE = 16'h8844;
		6206: SAMPLE = 16'h8776;
		6207: SAMPLE = 16'h86b3;
		6208: SAMPLE = 16'h85fc;
		6209: SAMPLE = 16'h854f;
		6210: SAMPLE = 16'h84ad;
		6211: SAMPLE = 16'h8416;
		6212: SAMPLE = 16'h838a;
		6213: SAMPLE = 16'h8308;
		6214: SAMPLE = 16'h8291;
		6215: SAMPLE = 16'h8224;
		6216: SAMPLE = 16'h81c1;
		6217: SAMPLE = 16'h8169;
		6218: SAMPLE = 16'h811b;
		6219: SAMPLE = 16'h80d6;
		6220: SAMPLE = 16'h809c;
		6221: SAMPLE = 16'h806b;
		6222: SAMPLE = 16'h8043;
		6223: SAMPLE = 16'h8025;
		6224: SAMPLE = 16'h800f;
		6225: SAMPLE = 16'h8003;
		6226: SAMPLE = 16'h8000;
		6227: SAMPLE = 16'h8004;
		6228: SAMPLE = 16'h8012;
		6229: SAMPLE = 16'h8027;
		6230: SAMPLE = 16'h8045;
		6231: SAMPLE = 16'h806a;
		6232: SAMPLE = 16'h8096;
		6233: SAMPLE = 16'h80ca;
		6234: SAMPLE = 16'h8106;
		6235: SAMPLE = 16'h8148;
		6236: SAMPLE = 16'h8190;
		6237: SAMPLE = 16'h81e0;
		6238: SAMPLE = 16'h8235;
		6239: SAMPLE = 16'h8290;
		6240: SAMPLE = 16'h82f1;
		6241: SAMPLE = 16'h8358;
		6242: SAMPLE = 16'h83c4;
		6243: SAMPLE = 16'h8435;
		6244: SAMPLE = 16'h84ab;
		6245: SAMPLE = 16'h8525;
		6246: SAMPLE = 16'h85a4;
		6247: SAMPLE = 16'h8627;
		6248: SAMPLE = 16'h86ad;
		6249: SAMPLE = 16'h8737;
		6250: SAMPLE = 16'h87c5;
		6251: SAMPLE = 16'h8855;
		6252: SAMPLE = 16'h88e9;
		6253: SAMPLE = 16'h897f;
		6254: SAMPLE = 16'h8a18;
		6255: SAMPLE = 16'h8ab2;
		6256: SAMPLE = 16'h8b4f;
		6257: SAMPLE = 16'h8bed;
		6258: SAMPLE = 16'h8c8d;
		6259: SAMPLE = 16'h8d2e;
		6260: SAMPLE = 16'h8dd0;
		6261: SAMPLE = 16'h8e73;
		6262: SAMPLE = 16'h8f16;
		6263: SAMPLE = 16'h8fba;
		6264: SAMPLE = 16'h905e;
		6265: SAMPLE = 16'h9102;
		6266: SAMPLE = 16'h91a5;
		6267: SAMPLE = 16'h9248;
		6268: SAMPLE = 16'h92ea;
		6269: SAMPLE = 16'h938c;
		6270: SAMPLE = 16'h942c;
		6271: SAMPLE = 16'h94cb;
		6272: SAMPLE = 16'h9568;
		6273: SAMPLE = 16'h9604;
		6274: SAMPLE = 16'h969e;
		6275: SAMPLE = 16'h9736;
		6276: SAMPLE = 16'h97cc;
		6277: SAMPLE = 16'h9860;
		6278: SAMPLE = 16'h98f1;
		6279: SAMPLE = 16'h9980;
		6280: SAMPLE = 16'h9a0b;
		6281: SAMPLE = 16'h9a94;
		6282: SAMPLE = 16'h9b1a;
		6283: SAMPLE = 16'h9b9d;
		6284: SAMPLE = 16'h9c1d;
		6285: SAMPLE = 16'h9c99;
		6286: SAMPLE = 16'h9d11;
		6287: SAMPLE = 16'h9d87;
		6288: SAMPLE = 16'h9df8;
		6289: SAMPLE = 16'h9e66;
		6290: SAMPLE = 16'h9ed0;
		6291: SAMPLE = 16'h9f36;
		6292: SAMPLE = 16'h9f98;
		6293: SAMPLE = 16'h9ff5;
		6294: SAMPLE = 16'ha04f;
		6295: SAMPLE = 16'ha0a5;
		6296: SAMPLE = 16'ha0f6;
		6297: SAMPLE = 16'ha143;
		6298: SAMPLE = 16'ha18c;
		6299: SAMPLE = 16'ha1d1;
		6300: SAMPLE = 16'ha211;
		6301: SAMPLE = 16'ha24d;
		6302: SAMPLE = 16'ha285;
		6303: SAMPLE = 16'ha2b8;
		6304: SAMPLE = 16'ha2e7;
		6305: SAMPLE = 16'ha311;
		6306: SAMPLE = 16'ha337;
		6307: SAMPLE = 16'ha359;
		6308: SAMPLE = 16'ha377;
		6309: SAMPLE = 16'ha390;
		6310: SAMPLE = 16'ha3a5;
		6311: SAMPLE = 16'ha3b6;
		6312: SAMPLE = 16'ha3c3;
		6313: SAMPLE = 16'ha3cb;
		6314: SAMPLE = 16'ha3d0;
		6315: SAMPLE = 16'ha3d1;
		6316: SAMPLE = 16'ha3cd;
		6317: SAMPLE = 16'ha3c6;
		6318: SAMPLE = 16'ha3bb;
		6319: SAMPLE = 16'ha3ad;
		6320: SAMPLE = 16'ha39b;
		6321: SAMPLE = 16'ha385;
		6322: SAMPLE = 16'ha36c;
		6323: SAMPLE = 16'ha350;
		6324: SAMPLE = 16'ha330;
		6325: SAMPLE = 16'ha30d;
		6326: SAMPLE = 16'ha2e7;
		6327: SAMPLE = 16'ha2bf;
		6328: SAMPLE = 16'ha293;
		6329: SAMPLE = 16'ha265;
		6330: SAMPLE = 16'ha234;
		6331: SAMPLE = 16'ha200;
		6332: SAMPLE = 16'ha1cb;
		6333: SAMPLE = 16'ha193;
		6334: SAMPLE = 16'ha159;
		6335: SAMPLE = 16'ha11c;
		6336: SAMPLE = 16'ha0df;
		6337: SAMPLE = 16'ha09f;
		6338: SAMPLE = 16'ha05d;
		6339: SAMPLE = 16'ha01b;
		6340: SAMPLE = 16'h9fd6;
		6341: SAMPLE = 16'h9f91;
		6342: SAMPLE = 16'h9f4b;
		6343: SAMPLE = 16'h9f03;
		6344: SAMPLE = 16'h9ebb;
		6345: SAMPLE = 16'h9e72;
		6346: SAMPLE = 16'h9e28;
		6347: SAMPLE = 16'h9dde;
		6348: SAMPLE = 16'h9d93;
		6349: SAMPLE = 16'h9d49;
		6350: SAMPLE = 16'h9cfe;
		6351: SAMPLE = 16'h9cb3;
		6352: SAMPLE = 16'h9c69;
		6353: SAMPLE = 16'h9c1f;
		6354: SAMPLE = 16'h9bd5;
		6355: SAMPLE = 16'h9b8c;
		6356: SAMPLE = 16'h9b43;
		6357: SAMPLE = 16'h9afc;
		6358: SAMPLE = 16'h9ab5;
		6359: SAMPLE = 16'h9a6f;
		6360: SAMPLE = 16'h9a2a;
		6361: SAMPLE = 16'h99e6;
		6362: SAMPLE = 16'h99a4;
		6363: SAMPLE = 16'h9963;
		6364: SAMPLE = 16'h9924;
		6365: SAMPLE = 16'h98e6;
		6366: SAMPLE = 16'h98aa;
		6367: SAMPLE = 16'h9870;
		6368: SAMPLE = 16'h9838;
		6369: SAMPLE = 16'h9801;
		6370: SAMPLE = 16'h97cd;
		6371: SAMPLE = 16'h979b;
		6372: SAMPLE = 16'h976b;
		6373: SAMPLE = 16'h973d;
		6374: SAMPLE = 16'h9711;
		6375: SAMPLE = 16'h96e8;
		6376: SAMPLE = 16'h96c2;
		6377: SAMPLE = 16'h969d;
		6378: SAMPLE = 16'h967c;
		6379: SAMPLE = 16'h965d;
		6380: SAMPLE = 16'h9640;
		6381: SAMPLE = 16'h9627;
		6382: SAMPLE = 16'h960f;
		6383: SAMPLE = 16'h95fb;
		6384: SAMPLE = 16'h95ea;
		6385: SAMPLE = 16'h95db;
		6386: SAMPLE = 16'h95cf;
		6387: SAMPLE = 16'h95c6;
		6388: SAMPLE = 16'h95bf;
		6389: SAMPLE = 16'h95bc;
		6390: SAMPLE = 16'h95bb;
		6391: SAMPLE = 16'h95bd;
		6392: SAMPLE = 16'h95c2;
		6393: SAMPLE = 16'h95ca;
		6394: SAMPLE = 16'h95d4;
		6395: SAMPLE = 16'h95e1;
		6396: SAMPLE = 16'h95f1;
		6397: SAMPLE = 16'h9604;
		6398: SAMPLE = 16'h961a;
		6399: SAMPLE = 16'h9632;
		6400: SAMPLE = 16'h964d;
		6401: SAMPLE = 16'h966a;
		6402: SAMPLE = 16'h968a;
		6403: SAMPLE = 16'h96ac;
		6404: SAMPLE = 16'h96d1;
		6405: SAMPLE = 16'h96f9;
		6406: SAMPLE = 16'h9722;
		6407: SAMPLE = 16'h974e;
		6408: SAMPLE = 16'h977d;
		6409: SAMPLE = 16'h97ad;
		6410: SAMPLE = 16'h97e0;
		6411: SAMPLE = 16'h9814;
		6412: SAMPLE = 16'h984b;
		6413: SAMPLE = 16'h9883;
		6414: SAMPLE = 16'h98be;
		6415: SAMPLE = 16'h98fa;
		6416: SAMPLE = 16'h9938;
		6417: SAMPLE = 16'h9977;
		6418: SAMPLE = 16'h99b8;
		6419: SAMPLE = 16'h99fa;
		6420: SAMPLE = 16'h9a3e;
		6421: SAMPLE = 16'h9a83;
		6422: SAMPLE = 16'h9ac9;
		6423: SAMPLE = 16'h9b11;
		6424: SAMPLE = 16'h9b59;
		6425: SAMPLE = 16'h9ba2;
		6426: SAMPLE = 16'h9bec;
		6427: SAMPLE = 16'h9c37;
		6428: SAMPLE = 16'h9c82;
		6429: SAMPLE = 16'h9cce;
		6430: SAMPLE = 16'h9d1b;
		6431: SAMPLE = 16'h9d68;
		6432: SAMPLE = 16'h9db5;
		6433: SAMPLE = 16'h9e02;
		6434: SAMPLE = 16'h9e4f;
		6435: SAMPLE = 16'h9e9d;
		6436: SAMPLE = 16'h9eea;
		6437: SAMPLE = 16'h9f37;
		6438: SAMPLE = 16'h9f84;
		6439: SAMPLE = 16'h9fd1;
		6440: SAMPLE = 16'ha01d;
		6441: SAMPLE = 16'ha069;
		6442: SAMPLE = 16'ha0b4;
		6443: SAMPLE = 16'ha0fe;
		6444: SAMPLE = 16'ha148;
		6445: SAMPLE = 16'ha191;
		6446: SAMPLE = 16'ha1d9;
		6447: SAMPLE = 16'ha220;
		6448: SAMPLE = 16'ha266;
		6449: SAMPLE = 16'ha2aa;
		6450: SAMPLE = 16'ha2ee;
		6451: SAMPLE = 16'ha330;
		6452: SAMPLE = 16'ha371;
		6453: SAMPLE = 16'ha3b1;
		6454: SAMPLE = 16'ha3ef;
		6455: SAMPLE = 16'ha42c;
		6456: SAMPLE = 16'ha467;
		6457: SAMPLE = 16'ha4a0;
		6458: SAMPLE = 16'ha4d8;
		6459: SAMPLE = 16'ha50e;
		6460: SAMPLE = 16'ha542;
		6461: SAMPLE = 16'ha574;
		6462: SAMPLE = 16'ha5a5;
		6463: SAMPLE = 16'ha5d4;
		6464: SAMPLE = 16'ha600;
		6465: SAMPLE = 16'ha62b;
		6466: SAMPLE = 16'ha654;
		6467: SAMPLE = 16'ha67b;
		6468: SAMPLE = 16'ha6a0;
		6469: SAMPLE = 16'ha6c2;
		6470: SAMPLE = 16'ha6e3;
		6471: SAMPLE = 16'ha701;
		6472: SAMPLE = 16'ha71e;
		6473: SAMPLE = 16'ha738;
		6474: SAMPLE = 16'ha751;
		6475: SAMPLE = 16'ha767;
		6476: SAMPLE = 16'ha77b;
		6477: SAMPLE = 16'ha78d;
		6478: SAMPLE = 16'ha79d;
		6479: SAMPLE = 16'ha7aa;
		6480: SAMPLE = 16'ha7b6;
		6481: SAMPLE = 16'ha7c0;
		6482: SAMPLE = 16'ha7c7;
		6483: SAMPLE = 16'ha7cd;
		6484: SAMPLE = 16'ha7d1;
		6485: SAMPLE = 16'ha7d2;
		6486: SAMPLE = 16'ha7d2;
		6487: SAMPLE = 16'ha7d0;
		6488: SAMPLE = 16'ha7cc;
		6489: SAMPLE = 16'ha7c6;
		6490: SAMPLE = 16'ha7be;
		6491: SAMPLE = 16'ha7b4;
		6492: SAMPLE = 16'ha7a9;
		6493: SAMPLE = 16'ha79c;
		6494: SAMPLE = 16'ha78e;
		6495: SAMPLE = 16'ha77e;
		6496: SAMPLE = 16'ha76c;
		6497: SAMPLE = 16'ha759;
		6498: SAMPLE = 16'ha744;
		6499: SAMPLE = 16'ha72f;
		6500: SAMPLE = 16'ha717;
		6501: SAMPLE = 16'ha6ff;
		6502: SAMPLE = 16'ha6e5;
		6503: SAMPLE = 16'ha6cb;
		6504: SAMPLE = 16'ha6af;
		6505: SAMPLE = 16'ha692;
		6506: SAMPLE = 16'ha674;
		6507: SAMPLE = 16'ha656;
		6508: SAMPLE = 16'ha637;
		6509: SAMPLE = 16'ha617;
		6510: SAMPLE = 16'ha5f6;
		6511: SAMPLE = 16'ha5d5;
		6512: SAMPLE = 16'ha5b3;
		6513: SAMPLE = 16'ha591;
		6514: SAMPLE = 16'ha56e;
		6515: SAMPLE = 16'ha54b;
		6516: SAMPLE = 16'ha528;
		6517: SAMPLE = 16'ha504;
		6518: SAMPLE = 16'ha4e1;
		6519: SAMPLE = 16'ha4be;
		6520: SAMPLE = 16'ha49a;
		6521: SAMPLE = 16'ha477;
		6522: SAMPLE = 16'ha454;
		6523: SAMPLE = 16'ha431;
		6524: SAMPLE = 16'ha40e;
		6525: SAMPLE = 16'ha3ec;
		6526: SAMPLE = 16'ha3cb;
		6527: SAMPLE = 16'ha3a9;
		6528: SAMPLE = 16'ha389;
		6529: SAMPLE = 16'ha369;
		6530: SAMPLE = 16'ha34a;
		6531: SAMPLE = 16'ha32b;
		6532: SAMPLE = 16'ha30e;
		6533: SAMPLE = 16'ha2f1;
		6534: SAMPLE = 16'ha2d5;
		6535: SAMPLE = 16'ha2ba;
		6536: SAMPLE = 16'ha2a0;
		6537: SAMPLE = 16'ha288;
		6538: SAMPLE = 16'ha270;
		6539: SAMPLE = 16'ha25a;
		6540: SAMPLE = 16'ha245;
		6541: SAMPLE = 16'ha231;
		6542: SAMPLE = 16'ha21e;
		6543: SAMPLE = 16'ha20d;
		6544: SAMPLE = 16'ha1fe;
		6545: SAMPLE = 16'ha1ef;
		6546: SAMPLE = 16'ha1e2;
		6547: SAMPLE = 16'ha1d7;
		6548: SAMPLE = 16'ha1cd;
		6549: SAMPLE = 16'ha1c5;
		6550: SAMPLE = 16'ha1be;
		6551: SAMPLE = 16'ha1b9;
		6552: SAMPLE = 16'ha1b6;
		6553: SAMPLE = 16'ha1b4;
		6554: SAMPLE = 16'ha1b4;
		6555: SAMPLE = 16'ha1b5;
		6556: SAMPLE = 16'ha1b9;
		6557: SAMPLE = 16'ha1bd;
		6558: SAMPLE = 16'ha1c4;
		6559: SAMPLE = 16'ha1cc;
		6560: SAMPLE = 16'ha1d6;
		6561: SAMPLE = 16'ha1e2;
		6562: SAMPLE = 16'ha1ef;
		6563: SAMPLE = 16'ha1fe;
		6564: SAMPLE = 16'ha20f;
		6565: SAMPLE = 16'ha221;
		6566: SAMPLE = 16'ha235;
		6567: SAMPLE = 16'ha24a;
		6568: SAMPLE = 16'ha261;
		6569: SAMPLE = 16'ha27a;
		6570: SAMPLE = 16'ha295;
		6571: SAMPLE = 16'ha2b0;
		6572: SAMPLE = 16'ha2ce;
		6573: SAMPLE = 16'ha2ed;
		6574: SAMPLE = 16'ha30d;
		6575: SAMPLE = 16'ha32f;
		6576: SAMPLE = 16'ha352;
		6577: SAMPLE = 16'ha376;
		6578: SAMPLE = 16'ha39c;
		6579: SAMPLE = 16'ha3c3;
		6580: SAMPLE = 16'ha3eb;
		6581: SAMPLE = 16'ha415;
		6582: SAMPLE = 16'ha43f;
		6583: SAMPLE = 16'ha46b;
		6584: SAMPLE = 16'ha498;
		6585: SAMPLE = 16'ha4c6;
		6586: SAMPLE = 16'ha4f5;
		6587: SAMPLE = 16'ha524;
		6588: SAMPLE = 16'ha555;
		6589: SAMPLE = 16'ha586;
		6590: SAMPLE = 16'ha5b8;
		6591: SAMPLE = 16'ha5eb;
		6592: SAMPLE = 16'ha61f;
		6593: SAMPLE = 16'ha653;
		6594: SAMPLE = 16'ha687;
		6595: SAMPLE = 16'ha6bc;
		6596: SAMPLE = 16'ha6f2;
		6597: SAMPLE = 16'ha728;
		6598: SAMPLE = 16'ha75e;
		6599: SAMPLE = 16'ha794;
		6600: SAMPLE = 16'ha7cb;
		6601: SAMPLE = 16'ha801;
		6602: SAMPLE = 16'ha838;
		6603: SAMPLE = 16'ha86f;
		6604: SAMPLE = 16'ha8a6;
		6605: SAMPLE = 16'ha8dc;
		6606: SAMPLE = 16'ha913;
		6607: SAMPLE = 16'ha949;
		6608: SAMPLE = 16'ha97f;
		6609: SAMPLE = 16'ha9b5;
		6610: SAMPLE = 16'ha9ea;
		6611: SAMPLE = 16'haa1f;
		6612: SAMPLE = 16'haa53;
		6613: SAMPLE = 16'haa87;
		6614: SAMPLE = 16'haabb;
		6615: SAMPLE = 16'haaed;
		6616: SAMPLE = 16'hab1f;
		6617: SAMPLE = 16'hab50;
		6618: SAMPLE = 16'hab81;
		6619: SAMPLE = 16'habb0;
		6620: SAMPLE = 16'habdf;
		6621: SAMPLE = 16'hac0d;
		6622: SAMPLE = 16'hac3a;
		6623: SAMPLE = 16'hac66;
		6624: SAMPLE = 16'hac91;
		6625: SAMPLE = 16'hacba;
		6626: SAMPLE = 16'hace3;
		6627: SAMPLE = 16'had0b;
		6628: SAMPLE = 16'had31;
		6629: SAMPLE = 16'had56;
		6630: SAMPLE = 16'had7a;
		6631: SAMPLE = 16'had9d;
		6632: SAMPLE = 16'hadbe;
		6633: SAMPLE = 16'hadde;
		6634: SAMPLE = 16'hadfd;
		6635: SAMPLE = 16'hae1b;
		6636: SAMPLE = 16'hae37;
		6637: SAMPLE = 16'hae52;
		6638: SAMPLE = 16'hae6b;
		6639: SAMPLE = 16'hae83;
		6640: SAMPLE = 16'hae9a;
		6641: SAMPLE = 16'haeaf;
		6642: SAMPLE = 16'haec3;
		6643: SAMPLE = 16'haed5;
		6644: SAMPLE = 16'haee6;
		6645: SAMPLE = 16'haef5;
		6646: SAMPLE = 16'haf04;
		6647: SAMPLE = 16'haf10;
		6648: SAMPLE = 16'haf1c;
		6649: SAMPLE = 16'haf26;
		6650: SAMPLE = 16'haf2e;
		6651: SAMPLE = 16'haf35;
		6652: SAMPLE = 16'haf3b;
		6653: SAMPLE = 16'haf40;
		6654: SAMPLE = 16'haf43;
		6655: SAMPLE = 16'haf45;
		6656: SAMPLE = 16'haf45;
		6657: SAMPLE = 16'haf45;
		6658: SAMPLE = 16'haf43;
		6659: SAMPLE = 16'haf40;
		6660: SAMPLE = 16'haf3c;
		6661: SAMPLE = 16'haf36;
		6662: SAMPLE = 16'haf30;
		6663: SAMPLE = 16'haf28;
		6664: SAMPLE = 16'haf20;
		6665: SAMPLE = 16'haf16;
		6666: SAMPLE = 16'haf0c;
		6667: SAMPLE = 16'haf00;
		6668: SAMPLE = 16'haef4;
		6669: SAMPLE = 16'haee7;
		6670: SAMPLE = 16'haed9;
		6671: SAMPLE = 16'haeca;
		6672: SAMPLE = 16'haeba;
		6673: SAMPLE = 16'haeaa;
		6674: SAMPLE = 16'hae99;
		6675: SAMPLE = 16'hae88;
		6676: SAMPLE = 16'hae76;
		6677: SAMPLE = 16'hae64;
		6678: SAMPLE = 16'hae51;
		6679: SAMPLE = 16'hae3d;
		6680: SAMPLE = 16'hae2a;
		6681: SAMPLE = 16'hae16;
		6682: SAMPLE = 16'hae02;
		6683: SAMPLE = 16'haded;
		6684: SAMPLE = 16'hadd9;
		6685: SAMPLE = 16'hadc4;
		6686: SAMPLE = 16'hadb0;
		6687: SAMPLE = 16'had9b;
		6688: SAMPLE = 16'had86;
		6689: SAMPLE = 16'had72;
		6690: SAMPLE = 16'had5d;
		6691: SAMPLE = 16'had49;
		6692: SAMPLE = 16'had35;
		6693: SAMPLE = 16'had21;
		6694: SAMPLE = 16'had0e;
		6695: SAMPLE = 16'hacfb;
		6696: SAMPLE = 16'hace8;
		6697: SAMPLE = 16'hacd6;
		6698: SAMPLE = 16'hacc5;
		6699: SAMPLE = 16'hacb4;
		6700: SAMPLE = 16'haca3;
		6701: SAMPLE = 16'hac93;
		6702: SAMPLE = 16'hac84;
		6703: SAMPLE = 16'hac76;
		6704: SAMPLE = 16'hac68;
		6705: SAMPLE = 16'hac5b;
		6706: SAMPLE = 16'hac4f;
		6707: SAMPLE = 16'hac44;
		6708: SAMPLE = 16'hac39;
		6709: SAMPLE = 16'hac30;
		6710: SAMPLE = 16'hac28;
		6711: SAMPLE = 16'hac20;
		6712: SAMPLE = 16'hac1a;
		6713: SAMPLE = 16'hac14;
		6714: SAMPLE = 16'hac10;
		6715: SAMPLE = 16'hac0d;
		6716: SAMPLE = 16'hac0a;
		6717: SAMPLE = 16'hac09;
		6718: SAMPLE = 16'hac09;
		6719: SAMPLE = 16'hac0b;
		6720: SAMPLE = 16'hac0d;
		6721: SAMPLE = 16'hac11;
		6722: SAMPLE = 16'hac15;
		6723: SAMPLE = 16'hac1b;
		6724: SAMPLE = 16'hac23;
		6725: SAMPLE = 16'hac2b;
		6726: SAMPLE = 16'hac35;
		6727: SAMPLE = 16'hac3f;
		6728: SAMPLE = 16'hac4b;
		6729: SAMPLE = 16'hac59;
		6730: SAMPLE = 16'hac67;
		6731: SAMPLE = 16'hac77;
		6732: SAMPLE = 16'hac88;
		6733: SAMPLE = 16'hac9a;
		6734: SAMPLE = 16'hacad;
		6735: SAMPLE = 16'hacc2;
		6736: SAMPLE = 16'hacd7;
		6737: SAMPLE = 16'hacee;
		6738: SAMPLE = 16'had06;
		6739: SAMPLE = 16'had1f;
		6740: SAMPLE = 16'had39;
		6741: SAMPLE = 16'had54;
		6742: SAMPLE = 16'had71;
		6743: SAMPLE = 16'had8e;
		6744: SAMPLE = 16'hadac;
		6745: SAMPLE = 16'hadcc;
		6746: SAMPLE = 16'hadec;
		6747: SAMPLE = 16'hae0d;
		6748: SAMPLE = 16'hae2f;
		6749: SAMPLE = 16'hae52;
		6750: SAMPLE = 16'hae76;
		6751: SAMPLE = 16'hae9a;
		6752: SAMPLE = 16'haec0;
		6753: SAMPLE = 16'haee6;
		6754: SAMPLE = 16'haf0d;
		6755: SAMPLE = 16'haf34;
		6756: SAMPLE = 16'haf5c;
		6757: SAMPLE = 16'haf85;
		6758: SAMPLE = 16'hafae;
		6759: SAMPLE = 16'hafd8;
		6760: SAMPLE = 16'hb002;
		6761: SAMPLE = 16'hb02c;
		6762: SAMPLE = 16'hb057;
		6763: SAMPLE = 16'hb082;
		6764: SAMPLE = 16'hb0ae;
		6765: SAMPLE = 16'hb0da;
		6766: SAMPLE = 16'hb106;
		6767: SAMPLE = 16'hb132;
		6768: SAMPLE = 16'hb15e;
		6769: SAMPLE = 16'hb18b;
		6770: SAMPLE = 16'hb1b7;
		6771: SAMPLE = 16'hb1e4;
		6772: SAMPLE = 16'hb210;
		6773: SAMPLE = 16'hb23c;
		6774: SAMPLE = 16'hb269;
		6775: SAMPLE = 16'hb295;
		6776: SAMPLE = 16'hb2c0;
		6777: SAMPLE = 16'hb2ec;
		6778: SAMPLE = 16'hb317;
		6779: SAMPLE = 16'hb342;
		6780: SAMPLE = 16'hb36c;
		6781: SAMPLE = 16'hb397;
		6782: SAMPLE = 16'hb3c0;
		6783: SAMPLE = 16'hb3e9;
		6784: SAMPLE = 16'hb412;
		6785: SAMPLE = 16'hb43a;
		6786: SAMPLE = 16'hb461;
		6787: SAMPLE = 16'hb488;
		6788: SAMPLE = 16'hb4ae;
		6789: SAMPLE = 16'hb4d4;
		6790: SAMPLE = 16'hb4f9;
		6791: SAMPLE = 16'hb51d;
		6792: SAMPLE = 16'hb540;
		6793: SAMPLE = 16'hb562;
		6794: SAMPLE = 16'hb584;
		6795: SAMPLE = 16'hb5a4;
		6796: SAMPLE = 16'hb5c4;
		6797: SAMPLE = 16'hb5e3;
		6798: SAMPLE = 16'hb601;
		6799: SAMPLE = 16'hb61e;
		6800: SAMPLE = 16'hb63a;
		6801: SAMPLE = 16'hb655;
		6802: SAMPLE = 16'hb66f;
		6803: SAMPLE = 16'hb687;
		6804: SAMPLE = 16'hb69f;
		6805: SAMPLE = 16'hb6b6;
		6806: SAMPLE = 16'hb6cc;
		6807: SAMPLE = 16'hb6e1;
		6808: SAMPLE = 16'hb6f4;
		6809: SAMPLE = 16'hb707;
		6810: SAMPLE = 16'hb719;
		6811: SAMPLE = 16'hb729;
		6812: SAMPLE = 16'hb738;
		6813: SAMPLE = 16'hb747;
		6814: SAMPLE = 16'hb754;
		6815: SAMPLE = 16'hb760;
		6816: SAMPLE = 16'hb76b;
		6817: SAMPLE = 16'hb775;
		6818: SAMPLE = 16'hb77e;
		6819: SAMPLE = 16'hb786;
		6820: SAMPLE = 16'hb78d;
		6821: SAMPLE = 16'hb793;
		6822: SAMPLE = 16'hb798;
		6823: SAMPLE = 16'hb79c;
		6824: SAMPLE = 16'hb79f;
		6825: SAMPLE = 16'hb7a1;
		6826: SAMPLE = 16'hb7a2;
		6827: SAMPLE = 16'hb7a2;
		6828: SAMPLE = 16'hb7a1;
		6829: SAMPLE = 16'hb7a0;
		6830: SAMPLE = 16'hb79d;
		6831: SAMPLE = 16'hb79a;
		6832: SAMPLE = 16'hb796;
		6833: SAMPLE = 16'hb791;
		6834: SAMPLE = 16'hb78c;
		6835: SAMPLE = 16'hb785;
		6836: SAMPLE = 16'hb77e;
		6837: SAMPLE = 16'hb777;
		6838: SAMPLE = 16'hb76f;
		6839: SAMPLE = 16'hb766;
		6840: SAMPLE = 16'hb75d;
		6841: SAMPLE = 16'hb753;
		6842: SAMPLE = 16'hb749;
		6843: SAMPLE = 16'hb73e;
		6844: SAMPLE = 16'hb733;
		6845: SAMPLE = 16'hb727;
		6846: SAMPLE = 16'hb71b;
		6847: SAMPLE = 16'hb70f;
		6848: SAMPLE = 16'hb703;
		6849: SAMPLE = 16'hb6f6;
		6850: SAMPLE = 16'hb6ea;
		6851: SAMPLE = 16'hb6dd;
		6852: SAMPLE = 16'hb6d0;
		6853: SAMPLE = 16'hb6c3;
		6854: SAMPLE = 16'hb6b6;
		6855: SAMPLE = 16'hb6a9;
		6856: SAMPLE = 16'hb69c;
		6857: SAMPLE = 16'hb68f;
		6858: SAMPLE = 16'hb682;
		6859: SAMPLE = 16'hb675;
		6860: SAMPLE = 16'hb669;
		6861: SAMPLE = 16'hb65d;
		6862: SAMPLE = 16'hb651;
		6863: SAMPLE = 16'hb645;
		6864: SAMPLE = 16'hb63a;
		6865: SAMPLE = 16'hb62f;
		6866: SAMPLE = 16'hb625;
		6867: SAMPLE = 16'hb61b;
		6868: SAMPLE = 16'hb611;
		6869: SAMPLE = 16'hb608;
		6870: SAMPLE = 16'hb600;
		6871: SAMPLE = 16'hb5f8;
		6872: SAMPLE = 16'hb5f1;
		6873: SAMPLE = 16'hb5ea;
		6874: SAMPLE = 16'hb5e4;
		6875: SAMPLE = 16'hb5df;
		6876: SAMPLE = 16'hb5da;
		6877: SAMPLE = 16'hb5d6;
		6878: SAMPLE = 16'hb5d3;
		6879: SAMPLE = 16'hb5d1;
		6880: SAMPLE = 16'hb5d0;
		6881: SAMPLE = 16'hb5cf;
		6882: SAMPLE = 16'hb5cf;
		6883: SAMPLE = 16'hb5d0;
		6884: SAMPLE = 16'hb5d2;
		6885: SAMPLE = 16'hb5d5;
		6886: SAMPLE = 16'hb5d9;
		6887: SAMPLE = 16'hb5dd;
		6888: SAMPLE = 16'hb5e3;
		6889: SAMPLE = 16'hb5e9;
		6890: SAMPLE = 16'hb5f1;
		6891: SAMPLE = 16'hb5f9;
		6892: SAMPLE = 16'hb603;
		6893: SAMPLE = 16'hb60d;
		6894: SAMPLE = 16'hb618;
		6895: SAMPLE = 16'hb625;
		6896: SAMPLE = 16'hb632;
		6897: SAMPLE = 16'hb640;
		6898: SAMPLE = 16'hb64f;
		6899: SAMPLE = 16'hb65f;
		6900: SAMPLE = 16'hb670;
		6901: SAMPLE = 16'hb682;
		6902: SAMPLE = 16'hb695;
		6903: SAMPLE = 16'hb6a9;
		6904: SAMPLE = 16'hb6be;
		6905: SAMPLE = 16'hb6d4;
		6906: SAMPLE = 16'hb6eb;
		6907: SAMPLE = 16'hb702;
		6908: SAMPLE = 16'hb71b;
		6909: SAMPLE = 16'hb734;
		6910: SAMPLE = 16'hb74e;
		6911: SAMPLE = 16'hb769;
		6912: SAMPLE = 16'hb785;
		6913: SAMPLE = 16'hb7a1;
		6914: SAMPLE = 16'hb7be;
		6915: SAMPLE = 16'hb7dc;
		6916: SAMPLE = 16'hb7fb;
		6917: SAMPLE = 16'hb81a;
		6918: SAMPLE = 16'hb83a;
		6919: SAMPLE = 16'hb85b;
		6920: SAMPLE = 16'hb87c;
		6921: SAMPLE = 16'hb89e;
		6922: SAMPLE = 16'hb8c0;
		6923: SAMPLE = 16'hb8e3;
		6924: SAMPLE = 16'hb907;
		6925: SAMPLE = 16'hb92a;
		6926: SAMPLE = 16'hb94f;
		6927: SAMPLE = 16'hb973;
		6928: SAMPLE = 16'hb998;
		6929: SAMPLE = 16'hb9bd;
		6930: SAMPLE = 16'hb9e3;
		6931: SAMPLE = 16'hba09;
		6932: SAMPLE = 16'hba2f;
		6933: SAMPLE = 16'hba55;
		6934: SAMPLE = 16'hba7b;
		6935: SAMPLE = 16'hbaa2;
		6936: SAMPLE = 16'hbac8;
		6937: SAMPLE = 16'hbaef;
		6938: SAMPLE = 16'hbb16;
		6939: SAMPLE = 16'hbb3c;
		6940: SAMPLE = 16'hbb63;
		6941: SAMPLE = 16'hbb89;
		6942: SAMPLE = 16'hbbb0;
		6943: SAMPLE = 16'hbbd6;
		6944: SAMPLE = 16'hbbfc;
		6945: SAMPLE = 16'hbc21;
		6946: SAMPLE = 16'hbc47;
		6947: SAMPLE = 16'hbc6c;
		6948: SAMPLE = 16'hbc91;
		6949: SAMPLE = 16'hbcb5;
		6950: SAMPLE = 16'hbcda;
		6951: SAMPLE = 16'hbcfd;
		6952: SAMPLE = 16'hbd21;
		6953: SAMPLE = 16'hbd43;
		6954: SAMPLE = 16'hbd66;
		6955: SAMPLE = 16'hbd87;
		6956: SAMPLE = 16'hbda9;
		6957: SAMPLE = 16'hbdc9;
		6958: SAMPLE = 16'hbde9;
		6959: SAMPLE = 16'hbe08;
		6960: SAMPLE = 16'hbe27;
		6961: SAMPLE = 16'hbe45;
		6962: SAMPLE = 16'hbe63;
		6963: SAMPLE = 16'hbe7f;
		6964: SAMPLE = 16'hbe9b;
		6965: SAMPLE = 16'hbeb6;
		6966: SAMPLE = 16'hbed1;
		6967: SAMPLE = 16'hbeea;
		6968: SAMPLE = 16'hbf03;
		6969: SAMPLE = 16'hbf1b;
		6970: SAMPLE = 16'hbf32;
		6971: SAMPLE = 16'hbf48;
		6972: SAMPLE = 16'hbf5e;
		6973: SAMPLE = 16'hbf72;
		6974: SAMPLE = 16'hbf86;
		6975: SAMPLE = 16'hbf99;
		6976: SAMPLE = 16'hbfab;
		6977: SAMPLE = 16'hbfbc;
		6978: SAMPLE = 16'hbfcc;
		6979: SAMPLE = 16'hbfdb;
		6980: SAMPLE = 16'hbfea;
		6981: SAMPLE = 16'hbff7;
		6982: SAMPLE = 16'hc004;
		6983: SAMPLE = 16'hc010;
		6984: SAMPLE = 16'hc01b;
		6985: SAMPLE = 16'hc025;
		6986: SAMPLE = 16'hc02e;
		6987: SAMPLE = 16'hc036;
		6988: SAMPLE = 16'hc03e;
		6989: SAMPLE = 16'hc044;
		6990: SAMPLE = 16'hc04a;
		6991: SAMPLE = 16'hc04f;
		6992: SAMPLE = 16'hc053;
		6993: SAMPLE = 16'hc057;
		6994: SAMPLE = 16'hc05a;
		6995: SAMPLE = 16'hc05c;
		6996: SAMPLE = 16'hc05d;
		6997: SAMPLE = 16'hc05d;
		6998: SAMPLE = 16'hc05d;
		6999: SAMPLE = 16'hc05d;
		7000: SAMPLE = 16'hc05b;
		7001: SAMPLE = 16'hc059;
		7002: SAMPLE = 16'hc057;
		7003: SAMPLE = 16'hc053;
		7004: SAMPLE = 16'hc050;
		7005: SAMPLE = 16'hc04b;
		7006: SAMPLE = 16'hc047;
		7007: SAMPLE = 16'hc042;
		7008: SAMPLE = 16'hc03c;
		7009: SAMPLE = 16'hc036;
		7010: SAMPLE = 16'hc02f;
		7011: SAMPLE = 16'hc029;
		7012: SAMPLE = 16'hc022;
		7013: SAMPLE = 16'hc01a;
		7014: SAMPLE = 16'hc013;
		7015: SAMPLE = 16'hc00b;
		7016: SAMPLE = 16'hc003;
		7017: SAMPLE = 16'hbffb;
		7018: SAMPLE = 16'hbff3;
		7019: SAMPLE = 16'hbfea;
		7020: SAMPLE = 16'hbfe2;
		7021: SAMPLE = 16'hbfd9;
		7022: SAMPLE = 16'hbfd1;
		7023: SAMPLE = 16'hbfc8;
		7024: SAMPLE = 16'hbfc0;
		7025: SAMPLE = 16'hbfb8;
		7026: SAMPLE = 16'hbfaf;
		7027: SAMPLE = 16'hbfa7;
		7028: SAMPLE = 16'hbfa0;
		7029: SAMPLE = 16'hbf98;
		7030: SAMPLE = 16'hbf91;
		7031: SAMPLE = 16'hbf89;
		7032: SAMPLE = 16'hbf83;
		7033: SAMPLE = 16'hbf7c;
		7034: SAMPLE = 16'hbf76;
		7035: SAMPLE = 16'hbf70;
		7036: SAMPLE = 16'hbf6b;
		7037: SAMPLE = 16'hbf66;
		7038: SAMPLE = 16'hbf62;
		7039: SAMPLE = 16'hbf5e;
		7040: SAMPLE = 16'hbf5b;
		7041: SAMPLE = 16'hbf58;
		7042: SAMPLE = 16'hbf56;
		7043: SAMPLE = 16'hbf54;
		7044: SAMPLE = 16'hbf53;
		7045: SAMPLE = 16'hbf53;
		7046: SAMPLE = 16'hbf53;
		7047: SAMPLE = 16'hbf54;
		7048: SAMPLE = 16'hbf55;
		7049: SAMPLE = 16'hbf58;
		7050: SAMPLE = 16'hbf5b;
		7051: SAMPLE = 16'hbf5f;
		7052: SAMPLE = 16'hbf63;
		7053: SAMPLE = 16'hbf68;
		7054: SAMPLE = 16'hbf6e;
		7055: SAMPLE = 16'hbf75;
		7056: SAMPLE = 16'hbf7d;
		7057: SAMPLE = 16'hbf85;
		7058: SAMPLE = 16'hbf8e;
		7059: SAMPLE = 16'hbf98;
		7060: SAMPLE = 16'hbfa3;
		7061: SAMPLE = 16'hbfaf;
		7062: SAMPLE = 16'hbfbb;
		7063: SAMPLE = 16'hbfc8;
		7064: SAMPLE = 16'hbfd6;
		7065: SAMPLE = 16'hbfe5;
		7066: SAMPLE = 16'hbff5;
		7067: SAMPLE = 16'hc005;
		7068: SAMPLE = 16'hc017;
		7069: SAMPLE = 16'hc029;
		7070: SAMPLE = 16'hc03b;
		7071: SAMPLE = 16'hc04f;
		7072: SAMPLE = 16'hc064;
		7073: SAMPLE = 16'hc079;
		7074: SAMPLE = 16'hc08f;
		7075: SAMPLE = 16'hc0a5;
		7076: SAMPLE = 16'hc0bd;
		7077: SAMPLE = 16'hc0d5;
		7078: SAMPLE = 16'hc0ee;
		7079: SAMPLE = 16'hc107;
		7080: SAMPLE = 16'hc121;
		7081: SAMPLE = 16'hc13c;
		7082: SAMPLE = 16'hc157;
		7083: SAMPLE = 16'hc173;
		7084: SAMPLE = 16'hc190;
		7085: SAMPLE = 16'hc1ad;
		7086: SAMPLE = 16'hc1cb;
		7087: SAMPLE = 16'hc1e9;
		7088: SAMPLE = 16'hc208;
		7089: SAMPLE = 16'hc227;
		7090: SAMPLE = 16'hc246;
		7091: SAMPLE = 16'hc266;
		7092: SAMPLE = 16'hc287;
		7093: SAMPLE = 16'hc2a8;
		7094: SAMPLE = 16'hc2c9;
		7095: SAMPLE = 16'hc2ea;
		7096: SAMPLE = 16'hc30c;
		7097: SAMPLE = 16'hc32e;
		7098: SAMPLE = 16'hc350;
		7099: SAMPLE = 16'hc372;
		7100: SAMPLE = 16'hc395;
		7101: SAMPLE = 16'hc3b8;
		7102: SAMPLE = 16'hc3db;
		7103: SAMPLE = 16'hc3fd;
		7104: SAMPLE = 16'hc420;
		7105: SAMPLE = 16'hc443;
		7106: SAMPLE = 16'hc466;
		7107: SAMPLE = 16'hc489;
		7108: SAMPLE = 16'hc4ac;
		7109: SAMPLE = 16'hc4cf;
		7110: SAMPLE = 16'hc4f1;
		7111: SAMPLE = 16'hc514;
		7112: SAMPLE = 16'hc536;
		7113: SAMPLE = 16'hc558;
		7114: SAMPLE = 16'hc57a;
		7115: SAMPLE = 16'hc59c;
		7116: SAMPLE = 16'hc5bd;
		7117: SAMPLE = 16'hc5de;
		7118: SAMPLE = 16'hc5fe;
		7119: SAMPLE = 16'hc61f;
		7120: SAMPLE = 16'hc63e;
		7121: SAMPLE = 16'hc65e;
		7122: SAMPLE = 16'hc67d;
		7123: SAMPLE = 16'hc69b;
		7124: SAMPLE = 16'hc6b9;
		7125: SAMPLE = 16'hc6d7;
		7126: SAMPLE = 16'hc6f4;
		7127: SAMPLE = 16'hc710;
		7128: SAMPLE = 16'hc72c;
		7129: SAMPLE = 16'hc747;
		7130: SAMPLE = 16'hc762;
		7131: SAMPLE = 16'hc77c;
		7132: SAMPLE = 16'hc795;
		7133: SAMPLE = 16'hc7ae;
		7134: SAMPLE = 16'hc7c6;
		7135: SAMPLE = 16'hc7dd;
		7136: SAMPLE = 16'hc7f4;
		7137: SAMPLE = 16'hc80a;
		7138: SAMPLE = 16'hc81f;
		7139: SAMPLE = 16'hc834;
		7140: SAMPLE = 16'hc848;
		7141: SAMPLE = 16'hc85b;
		7142: SAMPLE = 16'hc86d;
		7143: SAMPLE = 16'hc87e;
		7144: SAMPLE = 16'hc88f;
		7145: SAMPLE = 16'hc89f;
		7146: SAMPLE = 16'hc8ae;
		7147: SAMPLE = 16'hc8bd;
		7148: SAMPLE = 16'hc8cb;
		7149: SAMPLE = 16'hc8d8;
		7150: SAMPLE = 16'hc8e4;
		7151: SAMPLE = 16'hc8ef;
		7152: SAMPLE = 16'hc8fa;
		7153: SAMPLE = 16'hc904;
		7154: SAMPLE = 16'hc90d;
		7155: SAMPLE = 16'hc916;
		7156: SAMPLE = 16'hc91e;
		7157: SAMPLE = 16'hc925;
		7158: SAMPLE = 16'hc92b;
		7159: SAMPLE = 16'hc931;
		7160: SAMPLE = 16'hc936;
		7161: SAMPLE = 16'hc93b;
		7162: SAMPLE = 16'hc93e;
		7163: SAMPLE = 16'hc941;
		7164: SAMPLE = 16'hc944;
		7165: SAMPLE = 16'hc946;
		7166: SAMPLE = 16'hc947;
		7167: SAMPLE = 16'hc948;
		7168: SAMPLE = 16'hc948;
		7169: SAMPLE = 16'hc948;
		7170: SAMPLE = 16'hc947;
		7171: SAMPLE = 16'hc946;
		7172: SAMPLE = 16'hc944;
		7173: SAMPLE = 16'hc942;
		7174: SAMPLE = 16'hc940;
		7175: SAMPLE = 16'hc93d;
		7176: SAMPLE = 16'hc93a;
		7177: SAMPLE = 16'hc936;
		7178: SAMPLE = 16'hc932;
		7179: SAMPLE = 16'hc92e;
		7180: SAMPLE = 16'hc92a;
		7181: SAMPLE = 16'hc925;
		7182: SAMPLE = 16'hc920;
		7183: SAMPLE = 16'hc91b;
		7184: SAMPLE = 16'hc916;
		7185: SAMPLE = 16'hc911;
		7186: SAMPLE = 16'hc90b;
		7187: SAMPLE = 16'hc906;
		7188: SAMPLE = 16'hc900;
		7189: SAMPLE = 16'hc8fb;
		7190: SAMPLE = 16'hc8f5;
		7191: SAMPLE = 16'hc8f0;
		7192: SAMPLE = 16'hc8ea;
		7193: SAMPLE = 16'hc8e5;
		7194: SAMPLE = 16'hc8e0;
		7195: SAMPLE = 16'hc8db;
		7196: SAMPLE = 16'hc8d6;
		7197: SAMPLE = 16'hc8d1;
		7198: SAMPLE = 16'hc8cd;
		7199: SAMPLE = 16'hc8c9;
		7200: SAMPLE = 16'hc8c5;
		7201: SAMPLE = 16'hc8c2;
		7202: SAMPLE = 16'hc8be;
		7203: SAMPLE = 16'hc8bc;
		7204: SAMPLE = 16'hc8b9;
		7205: SAMPLE = 16'hc8b7;
		7206: SAMPLE = 16'hc8b5;
		7207: SAMPLE = 16'hc8b4;
		7208: SAMPLE = 16'hc8b4;
		7209: SAMPLE = 16'hc8b3;
		7210: SAMPLE = 16'hc8b4;
		7211: SAMPLE = 16'hc8b4;
		7212: SAMPLE = 16'hc8b6;
		7213: SAMPLE = 16'hc8b8;
		7214: SAMPLE = 16'hc8ba;
		7215: SAMPLE = 16'hc8bd;
		7216: SAMPLE = 16'hc8c1;
		7217: SAMPLE = 16'hc8c5;
		7218: SAMPLE = 16'hc8ca;
		7219: SAMPLE = 16'hc8d0;
		7220: SAMPLE = 16'hc8d6;
		7221: SAMPLE = 16'hc8dd;
		7222: SAMPLE = 16'hc8e4;
		7223: SAMPLE = 16'hc8ed;
		7224: SAMPLE = 16'hc8f6;
		7225: SAMPLE = 16'hc8ff;
		7226: SAMPLE = 16'hc90a;
		7227: SAMPLE = 16'hc915;
		7228: SAMPLE = 16'hc920;
		7229: SAMPLE = 16'hc92d;
		7230: SAMPLE = 16'hc93a;
		7231: SAMPLE = 16'hc948;
		7232: SAMPLE = 16'hc957;
		7233: SAMPLE = 16'hc966;
		7234: SAMPLE = 16'hc976;
		7235: SAMPLE = 16'hc987;
		7236: SAMPLE = 16'hc998;
		7237: SAMPLE = 16'hc9aa;
		7238: SAMPLE = 16'hc9bd;
		7239: SAMPLE = 16'hc9d1;
		7240: SAMPLE = 16'hc9e5;
		7241: SAMPLE = 16'hc9fa;
		7242: SAMPLE = 16'hca0f;
		7243: SAMPLE = 16'hca25;
		7244: SAMPLE = 16'hca3c;
		7245: SAMPLE = 16'hca54;
		7246: SAMPLE = 16'hca6c;
		7247: SAMPLE = 16'hca84;
		7248: SAMPLE = 16'hca9d;
		7249: SAMPLE = 16'hcab7;
		7250: SAMPLE = 16'hcad1;
		7251: SAMPLE = 16'hcaec;
		7252: SAMPLE = 16'hcb07;
		7253: SAMPLE = 16'hcb23;
		7254: SAMPLE = 16'hcb3f;
		7255: SAMPLE = 16'hcb5c;
		7256: SAMPLE = 16'hcb79;
		7257: SAMPLE = 16'hcb96;
		7258: SAMPLE = 16'hcbb4;
		7259: SAMPLE = 16'hcbd2;
		7260: SAMPLE = 16'hcbf1;
		7261: SAMPLE = 16'hcc0f;
		7262: SAMPLE = 16'hcc2e;
		7263: SAMPLE = 16'hcc4e;
		7264: SAMPLE = 16'hcc6d;
		7265: SAMPLE = 16'hcc8d;
		7266: SAMPLE = 16'hccad;
		7267: SAMPLE = 16'hcccd;
		7268: SAMPLE = 16'hcced;
		7269: SAMPLE = 16'hcd0e;
		7270: SAMPLE = 16'hcd2e;
		7271: SAMPLE = 16'hcd4f;
		7272: SAMPLE = 16'hcd6f;
		7273: SAMPLE = 16'hcd90;
		7274: SAMPLE = 16'hcdb0;
		7275: SAMPLE = 16'hcdd0;
		7276: SAMPLE = 16'hcdf1;
		7277: SAMPLE = 16'hce11;
		7278: SAMPLE = 16'hce31;
		7279: SAMPLE = 16'hce51;
		7280: SAMPLE = 16'hce71;
		7281: SAMPLE = 16'hce91;
		7282: SAMPLE = 16'hceb0;
		7283: SAMPLE = 16'hcecf;
		7284: SAMPLE = 16'hceee;
		7285: SAMPLE = 16'hcf0c;
		7286: SAMPLE = 16'hcf2b;
		7287: SAMPLE = 16'hcf48;
		7288: SAMPLE = 16'hcf66;
		7289: SAMPLE = 16'hcf83;
		7290: SAMPLE = 16'hcfa0;
		7291: SAMPLE = 16'hcfbc;
		7292: SAMPLE = 16'hcfd8;
		7293: SAMPLE = 16'hcff3;
		7294: SAMPLE = 16'hd00e;
		7295: SAMPLE = 16'hd028;
		7296: SAMPLE = 16'hd042;
		7297: SAMPLE = 16'hd05c;
		7298: SAMPLE = 16'hd074;
		7299: SAMPLE = 16'hd08c;
		7300: SAMPLE = 16'hd0a4;
		7301: SAMPLE = 16'hd0bb;
		7302: SAMPLE = 16'hd0d2;
		7303: SAMPLE = 16'hd0e7;
		7304: SAMPLE = 16'hd0fd;
		7305: SAMPLE = 16'hd111;
		7306: SAMPLE = 16'hd125;
		7307: SAMPLE = 16'hd138;
		7308: SAMPLE = 16'hd14b;
		7309: SAMPLE = 16'hd15d;
		7310: SAMPLE = 16'hd16e;
		7311: SAMPLE = 16'hd17f;
		7312: SAMPLE = 16'hd18f;
		7313: SAMPLE = 16'hd19e;
		7314: SAMPLE = 16'hd1ac;
		7315: SAMPLE = 16'hd1ba;
		7316: SAMPLE = 16'hd1c8;
		7317: SAMPLE = 16'hd1d4;
		7318: SAMPLE = 16'hd1e0;
		7319: SAMPLE = 16'hd1eb;
		7320: SAMPLE = 16'hd1f6;
		7321: SAMPLE = 16'hd200;
		7322: SAMPLE = 16'hd209;
		7323: SAMPLE = 16'hd212;
		7324: SAMPLE = 16'hd21a;
		7325: SAMPLE = 16'hd221;
		7326: SAMPLE = 16'hd228;
		7327: SAMPLE = 16'hd22e;
		7328: SAMPLE = 16'hd233;
		7329: SAMPLE = 16'hd238;
		7330: SAMPLE = 16'hd23d;
		7331: SAMPLE = 16'hd241;
		7332: SAMPLE = 16'hd244;
		7333: SAMPLE = 16'hd247;
		7334: SAMPLE = 16'hd249;
		7335: SAMPLE = 16'hd24b;
		7336: SAMPLE = 16'hd24c;
		7337: SAMPLE = 16'hd24d;
		7338: SAMPLE = 16'hd24e;
		7339: SAMPLE = 16'hd24e;
		7340: SAMPLE = 16'hd24d;
		7341: SAMPLE = 16'hd24d;
		7342: SAMPLE = 16'hd24c;
		7343: SAMPLE = 16'hd24a;
		7344: SAMPLE = 16'hd249;
		7345: SAMPLE = 16'hd247;
		7346: SAMPLE = 16'hd245;
		7347: SAMPLE = 16'hd242;
		7348: SAMPLE = 16'hd23f;
		7349: SAMPLE = 16'hd23d;
		7350: SAMPLE = 16'hd23a;
		7351: SAMPLE = 16'hd236;
		7352: SAMPLE = 16'hd233;
		7353: SAMPLE = 16'hd230;
		7354: SAMPLE = 16'hd22c;
		7355: SAMPLE = 16'hd229;
		7356: SAMPLE = 16'hd225;
		7357: SAMPLE = 16'hd222;
		7358: SAMPLE = 16'hd21e;
		7359: SAMPLE = 16'hd21b;
		7360: SAMPLE = 16'hd218;
		7361: SAMPLE = 16'hd215;
		7362: SAMPLE = 16'hd212;
		7363: SAMPLE = 16'hd20f;
		7364: SAMPLE = 16'hd20c;
		7365: SAMPLE = 16'hd209;
		7366: SAMPLE = 16'hd207;
		7367: SAMPLE = 16'hd205;
		7368: SAMPLE = 16'hd203;
		7369: SAMPLE = 16'hd202;
		7370: SAMPLE = 16'hd201;
		7371: SAMPLE = 16'hd200;
		7372: SAMPLE = 16'hd1ff;
		7373: SAMPLE = 16'hd1ff;
		7374: SAMPLE = 16'hd1ff;
		7375: SAMPLE = 16'hd200;
		7376: SAMPLE = 16'hd201;
		7377: SAMPLE = 16'hd203;
		7378: SAMPLE = 16'hd205;
		7379: SAMPLE = 16'hd207;
		7380: SAMPLE = 16'hd20a;
		7381: SAMPLE = 16'hd20e;
		7382: SAMPLE = 16'hd212;
		7383: SAMPLE = 16'hd217;
		7384: SAMPLE = 16'hd21c;
		7385: SAMPLE = 16'hd221;
		7386: SAMPLE = 16'hd228;
		7387: SAMPLE = 16'hd22f;
		7388: SAMPLE = 16'hd236;
		7389: SAMPLE = 16'hd23e;
		7390: SAMPLE = 16'hd247;
		7391: SAMPLE = 16'hd250;
		7392: SAMPLE = 16'hd25a;
		7393: SAMPLE = 16'hd265;
		7394: SAMPLE = 16'hd270;
		7395: SAMPLE = 16'hd27c;
		7396: SAMPLE = 16'hd289;
		7397: SAMPLE = 16'hd296;
		7398: SAMPLE = 16'hd2a4;
		7399: SAMPLE = 16'hd2b2;
		7400: SAMPLE = 16'hd2c1;
		7401: SAMPLE = 16'hd2d1;
		7402: SAMPLE = 16'hd2e1;
		7403: SAMPLE = 16'hd2f2;
		7404: SAMPLE = 16'hd304;
		7405: SAMPLE = 16'hd316;
		7406: SAMPLE = 16'hd329;
		7407: SAMPLE = 16'hd33c;
		7408: SAMPLE = 16'hd351;
		7409: SAMPLE = 16'hd365;
		7410: SAMPLE = 16'hd37a;
		7411: SAMPLE = 16'hd390;
		7412: SAMPLE = 16'hd3a7;
		7413: SAMPLE = 16'hd3be;
		7414: SAMPLE = 16'hd3d5;
		7415: SAMPLE = 16'hd3ed;
		7416: SAMPLE = 16'hd406;
		7417: SAMPLE = 16'hd41f;
		7418: SAMPLE = 16'hd438;
		7419: SAMPLE = 16'hd452;
		7420: SAMPLE = 16'hd46c;
		7421: SAMPLE = 16'hd487;
		7422: SAMPLE = 16'hd4a2;
		7423: SAMPLE = 16'hd4be;
		7424: SAMPLE = 16'hd4da;
		7425: SAMPLE = 16'hd4f6;
		7426: SAMPLE = 16'hd513;
		7427: SAMPLE = 16'hd52f;
		7428: SAMPLE = 16'hd54d;
		7429: SAMPLE = 16'hd56a;
		7430: SAMPLE = 16'hd588;
		7431: SAMPLE = 16'hd5a6;
		7432: SAMPLE = 16'hd5c4;
		7433: SAMPLE = 16'hd5e2;
		7434: SAMPLE = 16'hd600;
		7435: SAMPLE = 16'hd61f;
		7436: SAMPLE = 16'hd63e;
		7437: SAMPLE = 16'hd65c;
		7438: SAMPLE = 16'hd67b;
		7439: SAMPLE = 16'hd69a;
		7440: SAMPLE = 16'hd6b9;
		7441: SAMPLE = 16'hd6d8;
		7442: SAMPLE = 16'hd6f6;
		7443: SAMPLE = 16'hd715;
		7444: SAMPLE = 16'hd734;
		7445: SAMPLE = 16'hd752;
		7446: SAMPLE = 16'hd770;
		7447: SAMPLE = 16'hd78f;
		7448: SAMPLE = 16'hd7ad;
		7449: SAMPLE = 16'hd7cb;
		7450: SAMPLE = 16'hd7e8;
		7451: SAMPLE = 16'hd806;
		7452: SAMPLE = 16'hd823;
		7453: SAMPLE = 16'hd83f;
		7454: SAMPLE = 16'hd85c;
		7455: SAMPLE = 16'hd878;
		7456: SAMPLE = 16'hd894;
		7457: SAMPLE = 16'hd8af;
		7458: SAMPLE = 16'hd8ca;
		7459: SAMPLE = 16'hd8e5;
		7460: SAMPLE = 16'hd8ff;
		7461: SAMPLE = 16'hd919;
		7462: SAMPLE = 16'hd933;
		7463: SAMPLE = 16'hd94b;
		7464: SAMPLE = 16'hd964;
		7465: SAMPLE = 16'hd97c;
		7466: SAMPLE = 16'hd993;
		7467: SAMPLE = 16'hd9aa;
		7468: SAMPLE = 16'hd9c0;
		7469: SAMPLE = 16'hd9d6;
		7470: SAMPLE = 16'hd9eb;
		7471: SAMPLE = 16'hda00;
		7472: SAMPLE = 16'hda14;
		7473: SAMPLE = 16'hda28;
		7474: SAMPLE = 16'hda3b;
		7475: SAMPLE = 16'hda4d;
		7476: SAMPLE = 16'hda5f;
		7477: SAMPLE = 16'hda70;
		7478: SAMPLE = 16'hda80;
		7479: SAMPLE = 16'hda90;
		7480: SAMPLE = 16'hda9f;
		7481: SAMPLE = 16'hdaae;
		7482: SAMPLE = 16'hdabc;
		7483: SAMPLE = 16'hdaca;
		7484: SAMPLE = 16'hdad6;
		7485: SAMPLE = 16'hdae3;
		7486: SAMPLE = 16'hdaee;
		7487: SAMPLE = 16'hdaf9;
		7488: SAMPLE = 16'hdb03;
		7489: SAMPLE = 16'hdb0d;
		7490: SAMPLE = 16'hdb16;
		7491: SAMPLE = 16'hdb1f;
		7492: SAMPLE = 16'hdb27;
		7493: SAMPLE = 16'hdb2e;
		7494: SAMPLE = 16'hdb35;
		7495: SAMPLE = 16'hdb3c;
		7496: SAMPLE = 16'hdb42;
		7497: SAMPLE = 16'hdb47;
		7498: SAMPLE = 16'hdb4c;
		7499: SAMPLE = 16'hdb50;
		7500: SAMPLE = 16'hdb54;
		7501: SAMPLE = 16'hdb57;
		7502: SAMPLE = 16'hdb5a;
		7503: SAMPLE = 16'hdb5d;
		7504: SAMPLE = 16'hdb5f;
		7505: SAMPLE = 16'hdb60;
		7506: SAMPLE = 16'hdb62;
		7507: SAMPLE = 16'hdb63;
		7508: SAMPLE = 16'hdb63;
		7509: SAMPLE = 16'hdb63;
		7510: SAMPLE = 16'hdb63;
		7511: SAMPLE = 16'hdb63;
		7512: SAMPLE = 16'hdb62;
		7513: SAMPLE = 16'hdb62;
		7514: SAMPLE = 16'hdb61;
		7515: SAMPLE = 16'hdb5f;
		7516: SAMPLE = 16'hdb5e;
		7517: SAMPLE = 16'hdb5c;
		7518: SAMPLE = 16'hdb5b;
		7519: SAMPLE = 16'hdb59;
		7520: SAMPLE = 16'hdb57;
		7521: SAMPLE = 16'hdb55;
		7522: SAMPLE = 16'hdb53;
		7523: SAMPLE = 16'hdb51;
		7524: SAMPLE = 16'hdb4f;
		7525: SAMPLE = 16'hdb4c;
		7526: SAMPLE = 16'hdb4a;
		7527: SAMPLE = 16'hdb49;
		7528: SAMPLE = 16'hdb47;
		7529: SAMPLE = 16'hdb45;
		7530: SAMPLE = 16'hdb43;
		7531: SAMPLE = 16'hdb42;
		7532: SAMPLE = 16'hdb41;
		7533: SAMPLE = 16'hdb40;
		7534: SAMPLE = 16'hdb3f;
		7535: SAMPLE = 16'hdb3e;
		7536: SAMPLE = 16'hdb3e;
		7537: SAMPLE = 16'hdb3e;
		7538: SAMPLE = 16'hdb3e;
		7539: SAMPLE = 16'hdb3f;
		7540: SAMPLE = 16'hdb40;
		7541: SAMPLE = 16'hdb41;
		7542: SAMPLE = 16'hdb43;
		7543: SAMPLE = 16'hdb45;
		7544: SAMPLE = 16'hdb47;
		7545: SAMPLE = 16'hdb4a;
		7546: SAMPLE = 16'hdb4d;
		7547: SAMPLE = 16'hdb51;
		7548: SAMPLE = 16'hdb55;
		7549: SAMPLE = 16'hdb5a;
		7550: SAMPLE = 16'hdb5f;
		7551: SAMPLE = 16'hdb65;
		7552: SAMPLE = 16'hdb6b;
		7553: SAMPLE = 16'hdb72;
		7554: SAMPLE = 16'hdb7a;
		7555: SAMPLE = 16'hdb81;
		7556: SAMPLE = 16'hdb8a;
		7557: SAMPLE = 16'hdb93;
		7558: SAMPLE = 16'hdb9d;
		7559: SAMPLE = 16'hdba7;
		7560: SAMPLE = 16'hdbb1;
		7561: SAMPLE = 16'hdbbd;
		7562: SAMPLE = 16'hdbc9;
		7563: SAMPLE = 16'hdbd5;
		7564: SAMPLE = 16'hdbe2;
		7565: SAMPLE = 16'hdbf0;
		7566: SAMPLE = 16'hdbfe;
		7567: SAMPLE = 16'hdc0d;
		7568: SAMPLE = 16'hdc1d;
		7569: SAMPLE = 16'hdc2d;
		7570: SAMPLE = 16'hdc3e;
		7571: SAMPLE = 16'hdc4f;
		7572: SAMPLE = 16'hdc61;
		7573: SAMPLE = 16'hdc73;
		7574: SAMPLE = 16'hdc86;
		7575: SAMPLE = 16'hdc9a;
		7576: SAMPLE = 16'hdcae;
		7577: SAMPLE = 16'hdcc2;
		7578: SAMPLE = 16'hdcd8;
		7579: SAMPLE = 16'hdced;
		7580: SAMPLE = 16'hdd03;
		7581: SAMPLE = 16'hdd1a;
		7582: SAMPLE = 16'hdd31;
		7583: SAMPLE = 16'hdd49;
		7584: SAMPLE = 16'hdd61;
		7585: SAMPLE = 16'hdd7a;
		7586: SAMPLE = 16'hdd92;
		7587: SAMPLE = 16'hddac;
		7588: SAMPLE = 16'hddc6;
		7589: SAMPLE = 16'hdde0;
		7590: SAMPLE = 16'hddfa;
		7591: SAMPLE = 16'hde15;
		7592: SAMPLE = 16'hde30;
		7593: SAMPLE = 16'hde4c;
		7594: SAMPLE = 16'hde68;
		7595: SAMPLE = 16'hde84;
		7596: SAMPLE = 16'hdea0;
		7597: SAMPLE = 16'hdebd;
		7598: SAMPLE = 16'hded9;
		7599: SAMPLE = 16'hdef6;
		7600: SAMPLE = 16'hdf13;
		7601: SAMPLE = 16'hdf31;
		7602: SAMPLE = 16'hdf4e;
		7603: SAMPLE = 16'hdf6b;
		7604: SAMPLE = 16'hdf89;
		7605: SAMPLE = 16'hdfa7;
		7606: SAMPLE = 16'hdfc4;
		7607: SAMPLE = 16'hdfe2;
		7608: SAMPLE = 16'hdfff;
		7609: SAMPLE = 16'he01d;
		7610: SAMPLE = 16'he03b;
		7611: SAMPLE = 16'he058;
		7612: SAMPLE = 16'he076;
		7613: SAMPLE = 16'he093;
		7614: SAMPLE = 16'he0b0;
		7615: SAMPLE = 16'he0cd;
		7616: SAMPLE = 16'he0ea;
		7617: SAMPLE = 16'he106;
		7618: SAMPLE = 16'he123;
		7619: SAMPLE = 16'he13f;
		7620: SAMPLE = 16'he15b;
		7621: SAMPLE = 16'he176;
		7622: SAMPLE = 16'he191;
		7623: SAMPLE = 16'he1ac;
		7624: SAMPLE = 16'he1c7;
		7625: SAMPLE = 16'he1e1;
		7626: SAMPLE = 16'he1fb;
		7627: SAMPLE = 16'he215;
		7628: SAMPLE = 16'he22e;
		7629: SAMPLE = 16'he246;
		7630: SAMPLE = 16'he25f;
		7631: SAMPLE = 16'he276;
		7632: SAMPLE = 16'he28e;
		7633: SAMPLE = 16'he2a5;
		7634: SAMPLE = 16'he2bb;
		7635: SAMPLE = 16'he2d1;
		7636: SAMPLE = 16'he2e6;
		7637: SAMPLE = 16'he2fb;
		7638: SAMPLE = 16'he30f;
		7639: SAMPLE = 16'he323;
		7640: SAMPLE = 16'he337;
		7641: SAMPLE = 16'he349;
		7642: SAMPLE = 16'he35b;
		7643: SAMPLE = 16'he36d;
		7644: SAMPLE = 16'he37e;
		7645: SAMPLE = 16'he38e;
		7646: SAMPLE = 16'he39e;
		7647: SAMPLE = 16'he3ae;
		7648: SAMPLE = 16'he3bc;
		7649: SAMPLE = 16'he3ca;
		7650: SAMPLE = 16'he3d8;
		7651: SAMPLE = 16'he3e5;
		7652: SAMPLE = 16'he3f1;
		7653: SAMPLE = 16'he3fd;
		7654: SAMPLE = 16'he408;
		7655: SAMPLE = 16'he413;
		7656: SAMPLE = 16'he41d;
		7657: SAMPLE = 16'he427;
		7658: SAMPLE = 16'he430;
		7659: SAMPLE = 16'he439;
		7660: SAMPLE = 16'he440;
		7661: SAMPLE = 16'he448;
		7662: SAMPLE = 16'he44f;
		7663: SAMPLE = 16'he455;
		7664: SAMPLE = 16'he45b;
		7665: SAMPLE = 16'he461;
		7666: SAMPLE = 16'he466;
		7667: SAMPLE = 16'he46a;
		7668: SAMPLE = 16'he46e;
		7669: SAMPLE = 16'he472;
		7670: SAMPLE = 16'he475;
		7671: SAMPLE = 16'he478;
		7672: SAMPLE = 16'he47b;
		7673: SAMPLE = 16'he47d;
		7674: SAMPLE = 16'he47f;
		7675: SAMPLE = 16'he480;
		7676: SAMPLE = 16'he481;
		7677: SAMPLE = 16'he482;
		7678: SAMPLE = 16'he483;
		7679: SAMPLE = 16'he483;
		7680: SAMPLE = 16'he483;
		7681: SAMPLE = 16'he483;
		7682: SAMPLE = 16'he483;
		7683: SAMPLE = 16'he482;
		7684: SAMPLE = 16'he482;
		7685: SAMPLE = 16'he481;
		7686: SAMPLE = 16'he480;
		7687: SAMPLE = 16'he47f;
		7688: SAMPLE = 16'he47e;
		7689: SAMPLE = 16'he47d;
		7690: SAMPLE = 16'he47c;
		7691: SAMPLE = 16'he47b;
		7692: SAMPLE = 16'he47a;
		7693: SAMPLE = 16'he479;
		7694: SAMPLE = 16'he478;
		7695: SAMPLE = 16'he477;
		7696: SAMPLE = 16'he476;
		7697: SAMPLE = 16'he475;
		7698: SAMPLE = 16'he475;
		7699: SAMPLE = 16'he474;
		7700: SAMPLE = 16'he474;
		7701: SAMPLE = 16'he474;
		7702: SAMPLE = 16'he474;
		7703: SAMPLE = 16'he475;
		7704: SAMPLE = 16'he476;
		7705: SAMPLE = 16'he477;
		7706: SAMPLE = 16'he478;
		7707: SAMPLE = 16'he47a;
		7708: SAMPLE = 16'he47c;
		7709: SAMPLE = 16'he47e;
		7710: SAMPLE = 16'he481;
		7711: SAMPLE = 16'he484;
		7712: SAMPLE = 16'he487;
		7713: SAMPLE = 16'he48b;
		7714: SAMPLE = 16'he48f;
		7715: SAMPLE = 16'he494;
		7716: SAMPLE = 16'he499;
		7717: SAMPLE = 16'he49f;
		7718: SAMPLE = 16'he4a5;
		7719: SAMPLE = 16'he4ac;
		7720: SAMPLE = 16'he4b3;
		7721: SAMPLE = 16'he4ba;
		7722: SAMPLE = 16'he4c3;
		7723: SAMPLE = 16'he4cb;
		7724: SAMPLE = 16'he4d4;
		7725: SAMPLE = 16'he4de;
		7726: SAMPLE = 16'he4e9;
		7727: SAMPLE = 16'he4f3;
		7728: SAMPLE = 16'he4ff;
		7729: SAMPLE = 16'he50b;
		7730: SAMPLE = 16'he517;
		7731: SAMPLE = 16'he524;
		7732: SAMPLE = 16'he532;
		7733: SAMPLE = 16'he540;
		7734: SAMPLE = 16'he54f;
		7735: SAMPLE = 16'he55e;
		7736: SAMPLE = 16'he56e;
		7737: SAMPLE = 16'he57e;
		7738: SAMPLE = 16'he58f;
		7739: SAMPLE = 16'he5a1;
		7740: SAMPLE = 16'he5b3;
		7741: SAMPLE = 16'he5c6;
		7742: SAMPLE = 16'he5d9;
		7743: SAMPLE = 16'he5ec;
		7744: SAMPLE = 16'he601;
		7745: SAMPLE = 16'he615;
		7746: SAMPLE = 16'he62b;
		7747: SAMPLE = 16'he640;
		7748: SAMPLE = 16'he656;
		7749: SAMPLE = 16'he66d;
		7750: SAMPLE = 16'he684;
		7751: SAMPLE = 16'he69b;
		7752: SAMPLE = 16'he6b3;
		7753: SAMPLE = 16'he6cc;
		7754: SAMPLE = 16'he6e4;
		7755: SAMPLE = 16'he6fe;
		7756: SAMPLE = 16'he717;
		7757: SAMPLE = 16'he731;
		7758: SAMPLE = 16'he74b;
		7759: SAMPLE = 16'he765;
		7760: SAMPLE = 16'he780;
		7761: SAMPLE = 16'he79b;
		7762: SAMPLE = 16'he7b6;
		7763: SAMPLE = 16'he7d2;
		7764: SAMPLE = 16'he7ee;
		7765: SAMPLE = 16'he80a;
		7766: SAMPLE = 16'he826;
		7767: SAMPLE = 16'he842;
		7768: SAMPLE = 16'he85e;
		7769: SAMPLE = 16'he87b;
		7770: SAMPLE = 16'he898;
		7771: SAMPLE = 16'he8b4;
		7772: SAMPLE = 16'he8d1;
		7773: SAMPLE = 16'he8ee;
		7774: SAMPLE = 16'he90b;
		7775: SAMPLE = 16'he928;
		7776: SAMPLE = 16'he945;
		7777: SAMPLE = 16'he961;
		7778: SAMPLE = 16'he97e;
		7779: SAMPLE = 16'he99b;
		7780: SAMPLE = 16'he9b7;
		7781: SAMPLE = 16'he9d4;
		7782: SAMPLE = 16'he9f0;
		7783: SAMPLE = 16'hea0c;
		7784: SAMPLE = 16'hea28;
		7785: SAMPLE = 16'hea44;
		7786: SAMPLE = 16'hea5f;
		7787: SAMPLE = 16'hea7a;
		7788: SAMPLE = 16'hea95;
		7789: SAMPLE = 16'heab0;
		7790: SAMPLE = 16'heaca;
		7791: SAMPLE = 16'heae4;
		7792: SAMPLE = 16'heafe;
		7793: SAMPLE = 16'heb17;
		7794: SAMPLE = 16'heb30;
		7795: SAMPLE = 16'heb49;
		7796: SAMPLE = 16'heb61;
		7797: SAMPLE = 16'heb79;
		7798: SAMPLE = 16'heb91;
		7799: SAMPLE = 16'heba8;
		7800: SAMPLE = 16'hebbe;
		7801: SAMPLE = 16'hebd4;
		7802: SAMPLE = 16'hebea;
		7803: SAMPLE = 16'hebff;
		7804: SAMPLE = 16'hec13;
		7805: SAMPLE = 16'hec28;
		7806: SAMPLE = 16'hec3b;
		7807: SAMPLE = 16'hec4e;
		7808: SAMPLE = 16'hec61;
		7809: SAMPLE = 16'hec73;
		7810: SAMPLE = 16'hec84;
		7811: SAMPLE = 16'hec95;
		7812: SAMPLE = 16'heca6;
		7813: SAMPLE = 16'hecb6;
		7814: SAMPLE = 16'hecc5;
		7815: SAMPLE = 16'hecd4;
		7816: SAMPLE = 16'hece2;
		7817: SAMPLE = 16'hecf0;
		7818: SAMPLE = 16'hecfd;
		7819: SAMPLE = 16'hed0a;
		7820: SAMPLE = 16'hed16;
		7821: SAMPLE = 16'hed21;
		7822: SAMPLE = 16'hed2c;
		7823: SAMPLE = 16'hed36;
		7824: SAMPLE = 16'hed40;
		7825: SAMPLE = 16'hed4a;
		7826: SAMPLE = 16'hed53;
		7827: SAMPLE = 16'hed5b;
		7828: SAMPLE = 16'hed63;
		7829: SAMPLE = 16'hed6a;
		7830: SAMPLE = 16'hed71;
		7831: SAMPLE = 16'hed77;
		7832: SAMPLE = 16'hed7d;
		7833: SAMPLE = 16'hed83;
		7834: SAMPLE = 16'hed88;
		7835: SAMPLE = 16'hed8d;
		7836: SAMPLE = 16'hed91;
		7837: SAMPLE = 16'hed95;
		7838: SAMPLE = 16'hed98;
		7839: SAMPLE = 16'hed9b;
		7840: SAMPLE = 16'hed9e;
		7841: SAMPLE = 16'heda0;
		7842: SAMPLE = 16'heda2;
		7843: SAMPLE = 16'heda4;
		7844: SAMPLE = 16'heda6;
		7845: SAMPLE = 16'heda7;
		7846: SAMPLE = 16'heda8;
		7847: SAMPLE = 16'heda9;
		7848: SAMPLE = 16'heda9;
		7849: SAMPLE = 16'heda9;
		7850: SAMPLE = 16'hedaa;
		7851: SAMPLE = 16'hedaa;
		7852: SAMPLE = 16'heda9;
		7853: SAMPLE = 16'heda9;
		7854: SAMPLE = 16'heda9;
		7855: SAMPLE = 16'heda9;
		7856: SAMPLE = 16'heda8;
		7857: SAMPLE = 16'heda8;
		7858: SAMPLE = 16'heda7;
		7859: SAMPLE = 16'heda7;
		7860: SAMPLE = 16'heda6;
		7861: SAMPLE = 16'heda6;
		7862: SAMPLE = 16'heda6;
		7863: SAMPLE = 16'heda5;
		7864: SAMPLE = 16'heda5;
		7865: SAMPLE = 16'heda5;
		7866: SAMPLE = 16'heda5;
		7867: SAMPLE = 16'heda6;
		7868: SAMPLE = 16'heda6;
		7869: SAMPLE = 16'heda7;
		7870: SAMPLE = 16'heda8;
		7871: SAMPLE = 16'heda9;
		7872: SAMPLE = 16'hedab;
		7873: SAMPLE = 16'hedad;
		7874: SAMPLE = 16'hedaf;
		7875: SAMPLE = 16'hedb1;
		7876: SAMPLE = 16'hedb4;
		7877: SAMPLE = 16'hedb7;
		7878: SAMPLE = 16'hedba;
		7879: SAMPLE = 16'hedbe;
		7880: SAMPLE = 16'hedc2;
		7881: SAMPLE = 16'hedc7;
		7882: SAMPLE = 16'hedcc;
		7883: SAMPLE = 16'hedd1;
		7884: SAMPLE = 16'hedd7;
		7885: SAMPLE = 16'hedde;
		7886: SAMPLE = 16'hede4;
		7887: SAMPLE = 16'hedec;
		7888: SAMPLE = 16'hedf4;
		7889: SAMPLE = 16'hedfc;
		7890: SAMPLE = 16'hee05;
		7891: SAMPLE = 16'hee0e;
		7892: SAMPLE = 16'hee18;
		7893: SAMPLE = 16'hee22;
		7894: SAMPLE = 16'hee2d;
		7895: SAMPLE = 16'hee38;
		7896: SAMPLE = 16'hee44;
		7897: SAMPLE = 16'hee51;
		7898: SAMPLE = 16'hee5e;
		7899: SAMPLE = 16'hee6b;
		7900: SAMPLE = 16'hee79;
		7901: SAMPLE = 16'hee88;
		7902: SAMPLE = 16'hee97;
		7903: SAMPLE = 16'heea7;
		7904: SAMPLE = 16'heeb7;
		7905: SAMPLE = 16'heec8;
		7906: SAMPLE = 16'heed9;
		7907: SAMPLE = 16'heeeb;
		7908: SAMPLE = 16'heefd;
		7909: SAMPLE = 16'hef10;
		7910: SAMPLE = 16'hef24;
		7911: SAMPLE = 16'hef38;
		7912: SAMPLE = 16'hef4c;
		7913: SAMPLE = 16'hef61;
		7914: SAMPLE = 16'hef76;
		7915: SAMPLE = 16'hef8c;
		7916: SAMPLE = 16'hefa2;
		7917: SAMPLE = 16'hefb9;
		7918: SAMPLE = 16'hefd0;
		7919: SAMPLE = 16'hefe7;
		7920: SAMPLE = 16'hefff;
		7921: SAMPLE = 16'hf017;
		7922: SAMPLE = 16'hf030;
		7923: SAMPLE = 16'hf049;
		7924: SAMPLE = 16'hf062;
		7925: SAMPLE = 16'hf07c;
		7926: SAMPLE = 16'hf096;
		7927: SAMPLE = 16'hf0b0;
		7928: SAMPLE = 16'hf0cb;
		7929: SAMPLE = 16'hf0e6;
		7930: SAMPLE = 16'hf101;
		7931: SAMPLE = 16'hf11c;
		7932: SAMPLE = 16'hf137;
		7933: SAMPLE = 16'hf153;
		7934: SAMPLE = 16'hf16f;
		7935: SAMPLE = 16'hf18b;
		7936: SAMPLE = 16'hf1a7;
		7937: SAMPLE = 16'hf1c3;
		7938: SAMPLE = 16'hf1df;
		7939: SAMPLE = 16'hf1fb;
		7940: SAMPLE = 16'hf218;
		7941: SAMPLE = 16'hf234;
		7942: SAMPLE = 16'hf250;
		7943: SAMPLE = 16'hf26d;
		7944: SAMPLE = 16'hf289;
		7945: SAMPLE = 16'hf2a5;
		7946: SAMPLE = 16'hf2c1;
		7947: SAMPLE = 16'hf2dd;
		7948: SAMPLE = 16'hf2f9;
		7949: SAMPLE = 16'hf315;
		7950: SAMPLE = 16'hf331;
		7951: SAMPLE = 16'hf34c;
		7952: SAMPLE = 16'hf368;
		7953: SAMPLE = 16'hf383;
		7954: SAMPLE = 16'hf39e;
		7955: SAMPLE = 16'hf3b8;
		7956: SAMPLE = 16'hf3d3;
		7957: SAMPLE = 16'hf3ed;
		7958: SAMPLE = 16'hf406;
		7959: SAMPLE = 16'hf420;
		7960: SAMPLE = 16'hf439;
		7961: SAMPLE = 16'hf452;
		7962: SAMPLE = 16'hf46a;
		7963: SAMPLE = 16'hf482;
		7964: SAMPLE = 16'hf49a;
		7965: SAMPLE = 16'hf4b1;
		7966: SAMPLE = 16'hf4c8;
		7967: SAMPLE = 16'hf4de;
		7968: SAMPLE = 16'hf4f4;
		7969: SAMPLE = 16'hf509;
		7970: SAMPLE = 16'hf51e;
		7971: SAMPLE = 16'hf533;
		7972: SAMPLE = 16'hf547;
		7973: SAMPLE = 16'hf55a;
		7974: SAMPLE = 16'hf56d;
		7975: SAMPLE = 16'hf580;
		7976: SAMPLE = 16'hf592;
		7977: SAMPLE = 16'hf5a3;
		7978: SAMPLE = 16'hf5b4;
		7979: SAMPLE = 16'hf5c5;
		7980: SAMPLE = 16'hf5d5;
		7981: SAMPLE = 16'hf5e4;
		7982: SAMPLE = 16'hf5f3;
		7983: SAMPLE = 16'hf601;
		7984: SAMPLE = 16'hf60f;
		7985: SAMPLE = 16'hf61c;
		7986: SAMPLE = 16'hf629;
		7987: SAMPLE = 16'hf635;
		7988: SAMPLE = 16'hf641;
		7989: SAMPLE = 16'hf64c;
		7990: SAMPLE = 16'hf657;
		7991: SAMPLE = 16'hf661;
		7992: SAMPLE = 16'hf66b;
		7993: SAMPLE = 16'hf674;
		7994: SAMPLE = 16'hf67c;
		7995: SAMPLE = 16'hf684;
		7996: SAMPLE = 16'hf68c;
		7997: SAMPLE = 16'hf693;
		7998: SAMPLE = 16'hf69a;
		7999: SAMPLE = 16'hf6a0;
		8000: SAMPLE = 16'hf6a6;
		8001: SAMPLE = 16'hf6ab;
		8002: SAMPLE = 16'hf6b0;
		8003: SAMPLE = 16'hf6b5;
		8004: SAMPLE = 16'hf6b9;
		8005: SAMPLE = 16'hf6bd;
		8006: SAMPLE = 16'hf6c0;
		8007: SAMPLE = 16'hf6c3;
		8008: SAMPLE = 16'hf6c6;
		8009: SAMPLE = 16'hf6c8;
		8010: SAMPLE = 16'hf6cb;
		8011: SAMPLE = 16'hf6cc;
		8012: SAMPLE = 16'hf6ce;
		8013: SAMPLE = 16'hf6cf;
		8014: SAMPLE = 16'hf6d1;
		8015: SAMPLE = 16'hf6d1;
		8016: SAMPLE = 16'hf6d2;
		8017: SAMPLE = 16'hf6d3;
		8018: SAMPLE = 16'hf6d3;
		8019: SAMPLE = 16'hf6d3;
		8020: SAMPLE = 16'hf6d4;
		8021: SAMPLE = 16'hf6d4;
		8022: SAMPLE = 16'hf6d4;
		8023: SAMPLE = 16'hf6d4;
		8024: SAMPLE = 16'hf6d3;
		8025: SAMPLE = 16'hf6d3;
		8026: SAMPLE = 16'hf6d3;
		8027: SAMPLE = 16'hf6d3;
		8028: SAMPLE = 16'hf6d3;
		8029: SAMPLE = 16'hf6d3;
		8030: SAMPLE = 16'hf6d3;
		8031: SAMPLE = 16'hf6d3;
		8032: SAMPLE = 16'hf6d4;
		8033: SAMPLE = 16'hf6d4;
		8034: SAMPLE = 16'hf6d5;
		8035: SAMPLE = 16'hf6d6;
		8036: SAMPLE = 16'hf6d7;
		8037: SAMPLE = 16'hf6d8;
		8038: SAMPLE = 16'hf6da;
		8039: SAMPLE = 16'hf6db;
		8040: SAMPLE = 16'hf6dd;
		8041: SAMPLE = 16'hf6e0;
		8042: SAMPLE = 16'hf6e2;
		8043: SAMPLE = 16'hf6e5;
		8044: SAMPLE = 16'hf6e8;
		8045: SAMPLE = 16'hf6ec;
		8046: SAMPLE = 16'hf6f0;
		8047: SAMPLE = 16'hf6f4;
		8048: SAMPLE = 16'hf6f9;
		8049: SAMPLE = 16'hf6fe;
		8050: SAMPLE = 16'hf704;
		8051: SAMPLE = 16'hf70a;
		8052: SAMPLE = 16'hf710;
		8053: SAMPLE = 16'hf717;
		8054: SAMPLE = 16'hf71e;
		8055: SAMPLE = 16'hf726;
		8056: SAMPLE = 16'hf72f;
		8057: SAMPLE = 16'hf737;
		8058: SAMPLE = 16'hf741;
		8059: SAMPLE = 16'hf74b;
		8060: SAMPLE = 16'hf755;
		8061: SAMPLE = 16'hf760;
		8062: SAMPLE = 16'hf76b;
		8063: SAMPLE = 16'hf777;
		8064: SAMPLE = 16'hf783;
		8065: SAMPLE = 16'hf790;
		8066: SAMPLE = 16'hf79e;
		8067: SAMPLE = 16'hf7ac;
		8068: SAMPLE = 16'hf7ba;
		8069: SAMPLE = 16'hf7c9;
		8070: SAMPLE = 16'hf7d9;
		8071: SAMPLE = 16'hf7e9;
		8072: SAMPLE = 16'hf7fa;
		8073: SAMPLE = 16'hf80b;
		8074: SAMPLE = 16'hf81c;
		8075: SAMPLE = 16'hf82f;
		8076: SAMPLE = 16'hf841;
		8077: SAMPLE = 16'hf854;
		8078: SAMPLE = 16'hf868;
		8079: SAMPLE = 16'hf87c;
		8080: SAMPLE = 16'hf891;
		8081: SAMPLE = 16'hf8a6;
		8082: SAMPLE = 16'hf8bb;
		8083: SAMPLE = 16'hf8d1;
		8084: SAMPLE = 16'hf8e8;
		8085: SAMPLE = 16'hf8ff;
		8086: SAMPLE = 16'hf916;
		8087: SAMPLE = 16'hf92e;
		8088: SAMPLE = 16'hf946;
		8089: SAMPLE = 16'hf95e;
		8090: SAMPLE = 16'hf977;
		8091: SAMPLE = 16'hf990;
		8092: SAMPLE = 16'hf9a9;
		8093: SAMPLE = 16'hf9c3;
		8094: SAMPLE = 16'hf9dd;
		8095: SAMPLE = 16'hf9f7;
		8096: SAMPLE = 16'hfa12;
		8097: SAMPLE = 16'hfa2c;
		8098: SAMPLE = 16'hfa47;
		8099: SAMPLE = 16'hfa63;
		8100: SAMPLE = 16'hfa7e;
		8101: SAMPLE = 16'hfa99;
		8102: SAMPLE = 16'hfab5;
		8103: SAMPLE = 16'hfad1;
		8104: SAMPLE = 16'hfaed;
		8105: SAMPLE = 16'hfb09;
		8106: SAMPLE = 16'hfb25;
		8107: SAMPLE = 16'hfb41;
		8108: SAMPLE = 16'hfb5d;
		8109: SAMPLE = 16'hfb79;
		8110: SAMPLE = 16'hfb95;
		8111: SAMPLE = 16'hfbb1;
		8112: SAMPLE = 16'hfbcd;
		8113: SAMPLE = 16'hfbe9;
		8114: SAMPLE = 16'hfc05;
		8115: SAMPLE = 16'hfc21;
		8116: SAMPLE = 16'hfc3d;
		8117: SAMPLE = 16'hfc58;
		8118: SAMPLE = 16'hfc73;
		8119: SAMPLE = 16'hfc8e;
		8120: SAMPLE = 16'hfca9;
		8121: SAMPLE = 16'hfcc4;
		8122: SAMPLE = 16'hfcdf;
		8123: SAMPLE = 16'hfcf9;
		8124: SAMPLE = 16'hfd13;
		8125: SAMPLE = 16'hfd2c;
		8126: SAMPLE = 16'hfd46;
		8127: SAMPLE = 16'hfd5f;
		8128: SAMPLE = 16'hfd77;
		8129: SAMPLE = 16'hfd90;
		8130: SAMPLE = 16'hfda7;
		8131: SAMPLE = 16'hfdbf;
		8132: SAMPLE = 16'hfdd6;
		8133: SAMPLE = 16'hfded;
		8134: SAMPLE = 16'hfe03;
		8135: SAMPLE = 16'hfe19;
		8136: SAMPLE = 16'hfe2e;
		8137: SAMPLE = 16'hfe43;
		8138: SAMPLE = 16'hfe58;
		8139: SAMPLE = 16'hfe6c;
		8140: SAMPLE = 16'hfe80;
		8141: SAMPLE = 16'hfe93;
		8142: SAMPLE = 16'hfea5;
		8143: SAMPLE = 16'hfeb7;
		8144: SAMPLE = 16'hfec9;
		8145: SAMPLE = 16'hfeda;
		8146: SAMPLE = 16'hfeea;
		8147: SAMPLE = 16'hfefa;
		8148: SAMPLE = 16'hff0a;
		8149: SAMPLE = 16'hff19;
		8150: SAMPLE = 16'hff27;
		8151: SAMPLE = 16'hff35;
		8152: SAMPLE = 16'hff43;
		8153: SAMPLE = 16'hff4f;
		8154: SAMPLE = 16'hff5c;
		8155: SAMPLE = 16'hff67;
		8156: SAMPLE = 16'hff73;
		8157: SAMPLE = 16'hff7d;
		8158: SAMPLE = 16'hff88;
		8159: SAMPLE = 16'hff91;
		8160: SAMPLE = 16'hff9b;
		8161: SAMPLE = 16'hffa3;
		8162: SAMPLE = 16'hffac;
		8163: SAMPLE = 16'hffb4;
		8164: SAMPLE = 16'hffbb;
		8165: SAMPLE = 16'hffc2;
		8166: SAMPLE = 16'hffc8;
		8167: SAMPLE = 16'hffce;
		8168: SAMPLE = 16'hffd4;
		8169: SAMPLE = 16'hffd9;
		8170: SAMPLE = 16'hffdd;
		8171: SAMPLE = 16'hffe2;
		8172: SAMPLE = 16'hffe6;
		8173: SAMPLE = 16'hffe9;
		8174: SAMPLE = 16'hffed;
		8175: SAMPLE = 16'hfff0;
		8176: SAMPLE = 16'hfff2;
		8177: SAMPLE = 16'hfff5;
		8178: SAMPLE = 16'hfff7;
		8179: SAMPLE = 16'hfff8;
		8180: SAMPLE = 16'hfffa;
		8181: SAMPLE = 16'hfffb;
		8182: SAMPLE = 16'hfffc;
		8183: SAMPLE = 16'hfffd;
		8184: SAMPLE = 16'hfffe;
		8185: SAMPLE = 16'hfffe;
		8186: SAMPLE = 16'hffff;
		8187: SAMPLE = 16'hffff;
		8188: SAMPLE = 16'hffff;
		8189: SAMPLE = 16'hffff;
		8190: SAMPLE = 16'hffff;
		8191: SAMPLE = 16'hffff;
	endcase

end

endmodule
