// This is inefficient and should only be used in the testbench

module wave_table_test(
					  input logic [11:0] ADDR,
					  output logic [15:0] SAMPLE
					  );
					  
always_comb begin

	case(ADDR)
		0: SAMPLE = 16'h0;
		1: SAMPLE = 16'h32;
		2: SAMPLE = 16'h64;
		3: SAMPLE = 16'h96;
		4: SAMPLE = 16'hc9;
		5: SAMPLE = 16'hfb;
		6: SAMPLE = 16'h12d;
		7: SAMPLE = 16'h15f;
		8: SAMPLE = 16'h192;
		9: SAMPLE = 16'h1c4;
		10: SAMPLE = 16'h1f6;
		11: SAMPLE = 16'h228;
		12: SAMPLE = 16'h25b;
		13: SAMPLE = 16'h28d;
		14: SAMPLE = 16'h2bf;
		15: SAMPLE = 16'h2f1;
		16: SAMPLE = 16'h324;
		17: SAMPLE = 16'h356;
		18: SAMPLE = 16'h388;
		19: SAMPLE = 16'h3ba;
		20: SAMPLE = 16'h3ed;
		21: SAMPLE = 16'h41f;
		22: SAMPLE = 16'h451;
		23: SAMPLE = 16'h483;
		24: SAMPLE = 16'h4b6;
		25: SAMPLE = 16'h4e8;
		26: SAMPLE = 16'h51a;
		27: SAMPLE = 16'h54c;
		28: SAMPLE = 16'h57f;
		29: SAMPLE = 16'h5b1;
		30: SAMPLE = 16'h5e3;
		31: SAMPLE = 16'h615;
		32: SAMPLE = 16'h647;
		33: SAMPLE = 16'h67a;
		34: SAMPLE = 16'h6ac;
		35: SAMPLE = 16'h6de;
		36: SAMPLE = 16'h710;
		37: SAMPLE = 16'h742;
		38: SAMPLE = 16'h775;
		39: SAMPLE = 16'h7a7;
		40: SAMPLE = 16'h7d9;
		41: SAMPLE = 16'h80b;
		42: SAMPLE = 16'h83d;
		43: SAMPLE = 16'h86f;
		44: SAMPLE = 16'h8a2;
		45: SAMPLE = 16'h8d4;
		46: SAMPLE = 16'h906;
		47: SAMPLE = 16'h938;
		48: SAMPLE = 16'h96a;
		49: SAMPLE = 16'h99c;
		50: SAMPLE = 16'h9ce;
		51: SAMPLE = 16'ha00;
		52: SAMPLE = 16'ha33;
		53: SAMPLE = 16'ha65;
		54: SAMPLE = 16'ha97;
		55: SAMPLE = 16'hac9;
		56: SAMPLE = 16'hafb;
		57: SAMPLE = 16'hb2d;
		58: SAMPLE = 16'hb5f;
		59: SAMPLE = 16'hb91;
		60: SAMPLE = 16'hbc3;
		61: SAMPLE = 16'hbf5;
		62: SAMPLE = 16'hc27;
		63: SAMPLE = 16'hc59;
		64: SAMPLE = 16'hc8b;
		65: SAMPLE = 16'hcbd;
		66: SAMPLE = 16'hcef;
		67: SAMPLE = 16'hd21;
		68: SAMPLE = 16'hd53;
		69: SAMPLE = 16'hd85;
		70: SAMPLE = 16'hdb7;
		71: SAMPLE = 16'hde9;
		72: SAMPLE = 16'he1b;
		73: SAMPLE = 16'he4d;
		74: SAMPLE = 16'he7f;
		75: SAMPLE = 16'heb1;
		76: SAMPLE = 16'hee3;
		77: SAMPLE = 16'hf15;
		78: SAMPLE = 16'hf47;
		79: SAMPLE = 16'hf79;
		80: SAMPLE = 16'hfab;
		81: SAMPLE = 16'hfdd;
		82: SAMPLE = 16'h100e;
		83: SAMPLE = 16'h1040;
		84: SAMPLE = 16'h1072;
		85: SAMPLE = 16'h10a4;
		86: SAMPLE = 16'h10d6;
		87: SAMPLE = 16'h1108;
		88: SAMPLE = 16'h1139;
		89: SAMPLE = 16'h116b;
		90: SAMPLE = 16'h119d;
		91: SAMPLE = 16'h11cf;
		92: SAMPLE = 16'h1201;
		93: SAMPLE = 16'h1232;
		94: SAMPLE = 16'h1264;
		95: SAMPLE = 16'h1296;
		96: SAMPLE = 16'h12c8;
		97: SAMPLE = 16'h12f9;
		98: SAMPLE = 16'h132b;
		99: SAMPLE = 16'h135d;
		100: SAMPLE = 16'h138e;
		101: SAMPLE = 16'h13c0;
		102: SAMPLE = 16'h13f2;
		103: SAMPLE = 16'h1423;
		104: SAMPLE = 16'h1455;
		105: SAMPLE = 16'h1487;
		106: SAMPLE = 16'h14b8;
		107: SAMPLE = 16'h14ea;
		108: SAMPLE = 16'h151b;
		109: SAMPLE = 16'h154d;
		110: SAMPLE = 16'h157f;
		111: SAMPLE = 16'h15b0;
		112: SAMPLE = 16'h15e2;
		113: SAMPLE = 16'h1613;
		114: SAMPLE = 16'h1645;
		115: SAMPLE = 16'h1676;
		116: SAMPLE = 16'h16a8;
		117: SAMPLE = 16'h16d9;
		118: SAMPLE = 16'h170a;
		119: SAMPLE = 16'h173c;
		120: SAMPLE = 16'h176d;
		121: SAMPLE = 16'h179f;
		122: SAMPLE = 16'h17d0;
		123: SAMPLE = 16'h1802;
		124: SAMPLE = 16'h1833;
		125: SAMPLE = 16'h1864;
		126: SAMPLE = 16'h1896;
		127: SAMPLE = 16'h18c7;
		128: SAMPLE = 16'h18f8;
		129: SAMPLE = 16'h192a;
		130: SAMPLE = 16'h195b;
		131: SAMPLE = 16'h198c;
		132: SAMPLE = 16'h19bd;
		133: SAMPLE = 16'h19ef;
		134: SAMPLE = 16'h1a20;
		135: SAMPLE = 16'h1a51;
		136: SAMPLE = 16'h1a82;
		137: SAMPLE = 16'h1ab3;
		138: SAMPLE = 16'h1ae4;
		139: SAMPLE = 16'h1b16;
		140: SAMPLE = 16'h1b47;
		141: SAMPLE = 16'h1b78;
		142: SAMPLE = 16'h1ba9;
		143: SAMPLE = 16'h1bda;
		144: SAMPLE = 16'h1c0b;
		145: SAMPLE = 16'h1c3c;
		146: SAMPLE = 16'h1c6d;
		147: SAMPLE = 16'h1c9e;
		148: SAMPLE = 16'h1ccf;
		149: SAMPLE = 16'h1d00;
		150: SAMPLE = 16'h1d31;
		151: SAMPLE = 16'h1d62;
		152: SAMPLE = 16'h1d93;
		153: SAMPLE = 16'h1dc4;
		154: SAMPLE = 16'h1df5;
		155: SAMPLE = 16'h1e25;
		156: SAMPLE = 16'h1e56;
		157: SAMPLE = 16'h1e87;
		158: SAMPLE = 16'h1eb8;
		159: SAMPLE = 16'h1ee9;
		160: SAMPLE = 16'h1f19;
		161: SAMPLE = 16'h1f4a;
		162: SAMPLE = 16'h1f7b;
		163: SAMPLE = 16'h1fac;
		164: SAMPLE = 16'h1fdc;
		165: SAMPLE = 16'h200d;
		166: SAMPLE = 16'h203e;
		167: SAMPLE = 16'h206e;
		168: SAMPLE = 16'h209f;
		169: SAMPLE = 16'h20d0;
		170: SAMPLE = 16'h2100;
		171: SAMPLE = 16'h2131;
		172: SAMPLE = 16'h2161;
		173: SAMPLE = 16'h2192;
		174: SAMPLE = 16'h21c2;
		175: SAMPLE = 16'h21f3;
		176: SAMPLE = 16'h2223;
		177: SAMPLE = 16'h2254;
		178: SAMPLE = 16'h2284;
		179: SAMPLE = 16'h22b4;
		180: SAMPLE = 16'h22e5;
		181: SAMPLE = 16'h2315;
		182: SAMPLE = 16'h2345;
		183: SAMPLE = 16'h2376;
		184: SAMPLE = 16'h23a6;
		185: SAMPLE = 16'h23d6;
		186: SAMPLE = 16'h2407;
		187: SAMPLE = 16'h2437;
		188: SAMPLE = 16'h2467;
		189: SAMPLE = 16'h2497;
		190: SAMPLE = 16'h24c7;
		191: SAMPLE = 16'h24f7;
		192: SAMPLE = 16'h2528;
		193: SAMPLE = 16'h2558;
		194: SAMPLE = 16'h2588;
		195: SAMPLE = 16'h25b8;
		196: SAMPLE = 16'h25e8;
		197: SAMPLE = 16'h2618;
		198: SAMPLE = 16'h2648;
		199: SAMPLE = 16'h2678;
		200: SAMPLE = 16'h26a8;
		201: SAMPLE = 16'h26d8;
		202: SAMPLE = 16'h2707;
		203: SAMPLE = 16'h2737;
		204: SAMPLE = 16'h2767;
		205: SAMPLE = 16'h2797;
		206: SAMPLE = 16'h27c7;
		207: SAMPLE = 16'h27f6;
		208: SAMPLE = 16'h2826;
		209: SAMPLE = 16'h2856;
		210: SAMPLE = 16'h2886;
		211: SAMPLE = 16'h28b5;
		212: SAMPLE = 16'h28e5;
		213: SAMPLE = 16'h2915;
		214: SAMPLE = 16'h2944;
		215: SAMPLE = 16'h2974;
		216: SAMPLE = 16'h29a3;
		217: SAMPLE = 16'h29d3;
		218: SAMPLE = 16'h2a02;
		219: SAMPLE = 16'h2a32;
		220: SAMPLE = 16'h2a61;
		221: SAMPLE = 16'h2a91;
		222: SAMPLE = 16'h2ac0;
		223: SAMPLE = 16'h2aef;
		224: SAMPLE = 16'h2b1f;
		225: SAMPLE = 16'h2b4e;
		226: SAMPLE = 16'h2b7d;
		227: SAMPLE = 16'h2bad;
		228: SAMPLE = 16'h2bdc;
		229: SAMPLE = 16'h2c0b;
		230: SAMPLE = 16'h2c3a;
		231: SAMPLE = 16'h2c69;
		232: SAMPLE = 16'h2c98;
		233: SAMPLE = 16'h2cc8;
		234: SAMPLE = 16'h2cf7;
		235: SAMPLE = 16'h2d26;
		236: SAMPLE = 16'h2d55;
		237: SAMPLE = 16'h2d84;
		238: SAMPLE = 16'h2db3;
		239: SAMPLE = 16'h2de2;
		240: SAMPLE = 16'h2e11;
		241: SAMPLE = 16'h2e3f;
		242: SAMPLE = 16'h2e6e;
		243: SAMPLE = 16'h2e9d;
		244: SAMPLE = 16'h2ecc;
		245: SAMPLE = 16'h2efb;
		246: SAMPLE = 16'h2f29;
		247: SAMPLE = 16'h2f58;
		248: SAMPLE = 16'h2f87;
		249: SAMPLE = 16'h2fb5;
		250: SAMPLE = 16'h2fe4;
		251: SAMPLE = 16'h3013;
		252: SAMPLE = 16'h3041;
		253: SAMPLE = 16'h3070;
		254: SAMPLE = 16'h309e;
		255: SAMPLE = 16'h30cd;
		256: SAMPLE = 16'h30fb;
		257: SAMPLE = 16'h312a;
		258: SAMPLE = 16'h3158;
		259: SAMPLE = 16'h3186;
		260: SAMPLE = 16'h31b5;
		261: SAMPLE = 16'h31e3;
		262: SAMPLE = 16'h3211;
		263: SAMPLE = 16'h3240;
		264: SAMPLE = 16'h326e;
		265: SAMPLE = 16'h329c;
		266: SAMPLE = 16'h32ca;
		267: SAMPLE = 16'h32f8;
		268: SAMPLE = 16'h3326;
		269: SAMPLE = 16'h3354;
		270: SAMPLE = 16'h3382;
		271: SAMPLE = 16'h33b0;
		272: SAMPLE = 16'h33de;
		273: SAMPLE = 16'h340c;
		274: SAMPLE = 16'h343a;
		275: SAMPLE = 16'h3468;
		276: SAMPLE = 16'h3496;
		277: SAMPLE = 16'h34c4;
		278: SAMPLE = 16'h34f2;
		279: SAMPLE = 16'h351f;
		280: SAMPLE = 16'h354d;
		281: SAMPLE = 16'h357b;
		282: SAMPLE = 16'h35a8;
		283: SAMPLE = 16'h35d6;
		284: SAMPLE = 16'h3604;
		285: SAMPLE = 16'h3631;
		286: SAMPLE = 16'h365f;
		287: SAMPLE = 16'h368c;
		288: SAMPLE = 16'h36ba;
		289: SAMPLE = 16'h36e7;
		290: SAMPLE = 16'h3714;
		291: SAMPLE = 16'h3742;
		292: SAMPLE = 16'h376f;
		293: SAMPLE = 16'h379c;
		294: SAMPLE = 16'h37ca;
		295: SAMPLE = 16'h37f7;
		296: SAMPLE = 16'h3824;
		297: SAMPLE = 16'h3851;
		298: SAMPLE = 16'h387e;
		299: SAMPLE = 16'h38ab;
		300: SAMPLE = 16'h38d8;
		301: SAMPLE = 16'h3906;
		302: SAMPLE = 16'h3932;
		303: SAMPLE = 16'h395f;
		304: SAMPLE = 16'h398c;
		305: SAMPLE = 16'h39b9;
		306: SAMPLE = 16'h39e6;
		307: SAMPLE = 16'h3a13;
		308: SAMPLE = 16'h3a40;
		309: SAMPLE = 16'h3a6c;
		310: SAMPLE = 16'h3a99;
		311: SAMPLE = 16'h3ac6;
		312: SAMPLE = 16'h3af2;
		313: SAMPLE = 16'h3b1f;
		314: SAMPLE = 16'h3b4c;
		315: SAMPLE = 16'h3b78;
		316: SAMPLE = 16'h3ba5;
		317: SAMPLE = 16'h3bd1;
		318: SAMPLE = 16'h3bfd;
		319: SAMPLE = 16'h3c2a;
		320: SAMPLE = 16'h3c56;
		321: SAMPLE = 16'h3c83;
		322: SAMPLE = 16'h3caf;
		323: SAMPLE = 16'h3cdb;
		324: SAMPLE = 16'h3d07;
		325: SAMPLE = 16'h3d33;
		326: SAMPLE = 16'h3d60;
		327: SAMPLE = 16'h3d8c;
		328: SAMPLE = 16'h3db8;
		329: SAMPLE = 16'h3de4;
		330: SAMPLE = 16'h3e10;
		331: SAMPLE = 16'h3e3c;
		332: SAMPLE = 16'h3e68;
		333: SAMPLE = 16'h3e93;
		334: SAMPLE = 16'h3ebf;
		335: SAMPLE = 16'h3eeb;
		336: SAMPLE = 16'h3f17;
		337: SAMPLE = 16'h3f43;
		338: SAMPLE = 16'h3f6e;
		339: SAMPLE = 16'h3f9a;
		340: SAMPLE = 16'h3fc5;
		341: SAMPLE = 16'h3ff1;
		342: SAMPLE = 16'h401d;
		343: SAMPLE = 16'h4048;
		344: SAMPLE = 16'h4073;
		345: SAMPLE = 16'h409f;
		346: SAMPLE = 16'h40ca;
		347: SAMPLE = 16'h40f6;
		348: SAMPLE = 16'h4121;
		349: SAMPLE = 16'h414c;
		350: SAMPLE = 16'h4177;
		351: SAMPLE = 16'h41a2;
		352: SAMPLE = 16'h41ce;
		353: SAMPLE = 16'h41f9;
		354: SAMPLE = 16'h4224;
		355: SAMPLE = 16'h424f;
		356: SAMPLE = 16'h427a;
		357: SAMPLE = 16'h42a5;
		358: SAMPLE = 16'h42d0;
		359: SAMPLE = 16'h42fa;
		360: SAMPLE = 16'h4325;
		361: SAMPLE = 16'h4350;
		362: SAMPLE = 16'h437b;
		363: SAMPLE = 16'h43a5;
		364: SAMPLE = 16'h43d0;
		365: SAMPLE = 16'h43fb;
		366: SAMPLE = 16'h4425;
		367: SAMPLE = 16'h4450;
		368: SAMPLE = 16'h447a;
		369: SAMPLE = 16'h44a5;
		370: SAMPLE = 16'h44cf;
		371: SAMPLE = 16'h44fa;
		372: SAMPLE = 16'h4524;
		373: SAMPLE = 16'h454e;
		374: SAMPLE = 16'h4578;
		375: SAMPLE = 16'h45a3;
		376: SAMPLE = 16'h45cd;
		377: SAMPLE = 16'h45f7;
		378: SAMPLE = 16'h4621;
		379: SAMPLE = 16'h464b;
		380: SAMPLE = 16'h4675;
		381: SAMPLE = 16'h469f;
		382: SAMPLE = 16'h46c9;
		383: SAMPLE = 16'h46f3;
		384: SAMPLE = 16'h471c;
		385: SAMPLE = 16'h4746;
		386: SAMPLE = 16'h4770;
		387: SAMPLE = 16'h479a;
		388: SAMPLE = 16'h47c3;
		389: SAMPLE = 16'h47ed;
		390: SAMPLE = 16'h4816;
		391: SAMPLE = 16'h4840;
		392: SAMPLE = 16'h4869;
		393: SAMPLE = 16'h4893;
		394: SAMPLE = 16'h48bc;
		395: SAMPLE = 16'h48e6;
		396: SAMPLE = 16'h490f;
		397: SAMPLE = 16'h4938;
		398: SAMPLE = 16'h4961;
		399: SAMPLE = 16'h498a;
		400: SAMPLE = 16'h49b4;
		401: SAMPLE = 16'h49dd;
		402: SAMPLE = 16'h4a06;
		403: SAMPLE = 16'h4a2f;
		404: SAMPLE = 16'h4a58;
		405: SAMPLE = 16'h4a81;
		406: SAMPLE = 16'h4aa9;
		407: SAMPLE = 16'h4ad2;
		408: SAMPLE = 16'h4afb;
		409: SAMPLE = 16'h4b24;
		410: SAMPLE = 16'h4b4c;
		411: SAMPLE = 16'h4b75;
		412: SAMPLE = 16'h4b9e;
		413: SAMPLE = 16'h4bc6;
		414: SAMPLE = 16'h4bef;
		415: SAMPLE = 16'h4c17;
		416: SAMPLE = 16'h4c3f;
		417: SAMPLE = 16'h4c68;
		418: SAMPLE = 16'h4c90;
		419: SAMPLE = 16'h4cb8;
		420: SAMPLE = 16'h4ce1;
		421: SAMPLE = 16'h4d09;
		422: SAMPLE = 16'h4d31;
		423: SAMPLE = 16'h4d59;
		424: SAMPLE = 16'h4d81;
		425: SAMPLE = 16'h4da9;
		426: SAMPLE = 16'h4dd1;
		427: SAMPLE = 16'h4df9;
		428: SAMPLE = 16'h4e21;
		429: SAMPLE = 16'h4e48;
		430: SAMPLE = 16'h4e70;
		431: SAMPLE = 16'h4e98;
		432: SAMPLE = 16'h4ebf;
		433: SAMPLE = 16'h4ee7;
		434: SAMPLE = 16'h4f0f;
		435: SAMPLE = 16'h4f36;
		436: SAMPLE = 16'h4f5e;
		437: SAMPLE = 16'h4f85;
		438: SAMPLE = 16'h4fac;
		439: SAMPLE = 16'h4fd4;
		440: SAMPLE = 16'h4ffb;
		441: SAMPLE = 16'h5022;
		442: SAMPLE = 16'h5049;
		443: SAMPLE = 16'h5070;
		444: SAMPLE = 16'h5097;
		445: SAMPLE = 16'h50bf;
		446: SAMPLE = 16'h50e5;
		447: SAMPLE = 16'h510c;
		448: SAMPLE = 16'h5133;
		449: SAMPLE = 16'h515a;
		450: SAMPLE = 16'h5181;
		451: SAMPLE = 16'h51a8;
		452: SAMPLE = 16'h51ce;
		453: SAMPLE = 16'h51f5;
		454: SAMPLE = 16'h521c;
		455: SAMPLE = 16'h5242;
		456: SAMPLE = 16'h5269;
		457: SAMPLE = 16'h528f;
		458: SAMPLE = 16'h52b5;
		459: SAMPLE = 16'h52dc;
		460: SAMPLE = 16'h5302;
		461: SAMPLE = 16'h5328;
		462: SAMPLE = 16'h534e;
		463: SAMPLE = 16'h5375;
		464: SAMPLE = 16'h539b;
		465: SAMPLE = 16'h53c1;
		466: SAMPLE = 16'h53e7;
		467: SAMPLE = 16'h540d;
		468: SAMPLE = 16'h5433;
		469: SAMPLE = 16'h5458;
		470: SAMPLE = 16'h547e;
		471: SAMPLE = 16'h54a4;
		472: SAMPLE = 16'h54ca;
		473: SAMPLE = 16'h54ef;
		474: SAMPLE = 16'h5515;
		475: SAMPLE = 16'h553a;
		476: SAMPLE = 16'h5560;
		477: SAMPLE = 16'h5585;
		478: SAMPLE = 16'h55ab;
		479: SAMPLE = 16'h55d0;
		480: SAMPLE = 16'h55f5;
		481: SAMPLE = 16'h561a;
		482: SAMPLE = 16'h5640;
		483: SAMPLE = 16'h5665;
		484: SAMPLE = 16'h568a;
		485: SAMPLE = 16'h56af;
		486: SAMPLE = 16'h56d4;
		487: SAMPLE = 16'h56f9;
		488: SAMPLE = 16'h571d;
		489: SAMPLE = 16'h5742;
		490: SAMPLE = 16'h5767;
		491: SAMPLE = 16'h578c;
		492: SAMPLE = 16'h57b0;
		493: SAMPLE = 16'h57d5;
		494: SAMPLE = 16'h57f9;
		495: SAMPLE = 16'h581e;
		496: SAMPLE = 16'h5842;
		497: SAMPLE = 16'h5867;
		498: SAMPLE = 16'h588b;
		499: SAMPLE = 16'h58af;
		500: SAMPLE = 16'h58d4;
		501: SAMPLE = 16'h58f8;
		502: SAMPLE = 16'h591c;
		503: SAMPLE = 16'h5940;
		504: SAMPLE = 16'h5964;
		505: SAMPLE = 16'h5988;
		506: SAMPLE = 16'h59ac;
		507: SAMPLE = 16'h59d0;
		508: SAMPLE = 16'h59f3;
		509: SAMPLE = 16'h5a17;
		510: SAMPLE = 16'h5a3b;
		511: SAMPLE = 16'h5a5e;
		512: SAMPLE = 16'h5a82;
		513: SAMPLE = 16'h5aa5;
		514: SAMPLE = 16'h5ac9;
		515: SAMPLE = 16'h5aec;
		516: SAMPLE = 16'h5b10;
		517: SAMPLE = 16'h5b33;
		518: SAMPLE = 16'h5b56;
		519: SAMPLE = 16'h5b79;
		520: SAMPLE = 16'h5b9d;
		521: SAMPLE = 16'h5bc0;
		522: SAMPLE = 16'h5be3;
		523: SAMPLE = 16'h5c06;
		524: SAMPLE = 16'h5c29;
		525: SAMPLE = 16'h5c4b;
		526: SAMPLE = 16'h5c6e;
		527: SAMPLE = 16'h5c91;
		528: SAMPLE = 16'h5cb4;
		529: SAMPLE = 16'h5cd6;
		530: SAMPLE = 16'h5cf9;
		531: SAMPLE = 16'h5d1b;
		532: SAMPLE = 16'h5d3e;
		533: SAMPLE = 16'h5d60;
		534: SAMPLE = 16'h5d83;
		535: SAMPLE = 16'h5da5;
		536: SAMPLE = 16'h5dc7;
		537: SAMPLE = 16'h5de9;
		538: SAMPLE = 16'h5e0b;
		539: SAMPLE = 16'h5e2d;
		540: SAMPLE = 16'h5e50;
		541: SAMPLE = 16'h5e71;
		542: SAMPLE = 16'h5e93;
		543: SAMPLE = 16'h5eb5;
		544: SAMPLE = 16'h5ed7;
		545: SAMPLE = 16'h5ef9;
		546: SAMPLE = 16'h5f1a;
		547: SAMPLE = 16'h5f3c;
		548: SAMPLE = 16'h5f5e;
		549: SAMPLE = 16'h5f7f;
		550: SAMPLE = 16'h5fa0;
		551: SAMPLE = 16'h5fc2;
		552: SAMPLE = 16'h5fe3;
		553: SAMPLE = 16'h6004;
		554: SAMPLE = 16'h6026;
		555: SAMPLE = 16'h6047;
		556: SAMPLE = 16'h6068;
		557: SAMPLE = 16'h6089;
		558: SAMPLE = 16'h60aa;
		559: SAMPLE = 16'h60cb;
		560: SAMPLE = 16'h60ec;
		561: SAMPLE = 16'h610d;
		562: SAMPLE = 16'h612d;
		563: SAMPLE = 16'h614e;
		564: SAMPLE = 16'h616f;
		565: SAMPLE = 16'h618f;
		566: SAMPLE = 16'h61b0;
		567: SAMPLE = 16'h61d0;
		568: SAMPLE = 16'h61f1;
		569: SAMPLE = 16'h6211;
		570: SAMPLE = 16'h6231;
		571: SAMPLE = 16'h6251;
		572: SAMPLE = 16'h6271;
		573: SAMPLE = 16'h6292;
		574: SAMPLE = 16'h62b2;
		575: SAMPLE = 16'h62d2;
		576: SAMPLE = 16'h62f2;
		577: SAMPLE = 16'h6311;
		578: SAMPLE = 16'h6331;
		579: SAMPLE = 16'h6351;
		580: SAMPLE = 16'h6371;
		581: SAMPLE = 16'h6390;
		582: SAMPLE = 16'h63b0;
		583: SAMPLE = 16'h63cf;
		584: SAMPLE = 16'h63ef;
		585: SAMPLE = 16'h640e;
		586: SAMPLE = 16'h642d;
		587: SAMPLE = 16'h644d;
		588: SAMPLE = 16'h646c;
		589: SAMPLE = 16'h648b;
		590: SAMPLE = 16'h64aa;
		591: SAMPLE = 16'h64c9;
		592: SAMPLE = 16'h64e8;
		593: SAMPLE = 16'h6507;
		594: SAMPLE = 16'h6526;
		595: SAMPLE = 16'h6545;
		596: SAMPLE = 16'h6563;
		597: SAMPLE = 16'h6582;
		598: SAMPLE = 16'h65a0;
		599: SAMPLE = 16'h65bf;
		600: SAMPLE = 16'h65dd;
		601: SAMPLE = 16'h65fc;
		602: SAMPLE = 16'h661a;
		603: SAMPLE = 16'h6639;
		604: SAMPLE = 16'h6657;
		605: SAMPLE = 16'h6675;
		606: SAMPLE = 16'h6693;
		607: SAMPLE = 16'h66b1;
		608: SAMPLE = 16'h66cf;
		609: SAMPLE = 16'h66ed;
		610: SAMPLE = 16'h670b;
		611: SAMPLE = 16'h6729;
		612: SAMPLE = 16'h6746;
		613: SAMPLE = 16'h6764;
		614: SAMPLE = 16'h6782;
		615: SAMPLE = 16'h679f;
		616: SAMPLE = 16'h67bd;
		617: SAMPLE = 16'h67da;
		618: SAMPLE = 16'h67f7;
		619: SAMPLE = 16'h6815;
		620: SAMPLE = 16'h6832;
		621: SAMPLE = 16'h684f;
		622: SAMPLE = 16'h686c;
		623: SAMPLE = 16'h6889;
		624: SAMPLE = 16'h68a6;
		625: SAMPLE = 16'h68c3;
		626: SAMPLE = 16'h68e0;
		627: SAMPLE = 16'h68fd;
		628: SAMPLE = 16'h6919;
		629: SAMPLE = 16'h6936;
		630: SAMPLE = 16'h6953;
		631: SAMPLE = 16'h696f;
		632: SAMPLE = 16'h698c;
		633: SAMPLE = 16'h69a8;
		634: SAMPLE = 16'h69c4;
		635: SAMPLE = 16'h69e1;
		636: SAMPLE = 16'h69fd;
		637: SAMPLE = 16'h6a19;
		638: SAMPLE = 16'h6a35;
		639: SAMPLE = 16'h6a51;
		640: SAMPLE = 16'h6a6d;
		641: SAMPLE = 16'h6a89;
		642: SAMPLE = 16'h6aa5;
		643: SAMPLE = 16'h6ac1;
		644: SAMPLE = 16'h6adc;
		645: SAMPLE = 16'h6af8;
		646: SAMPLE = 16'h6b13;
		647: SAMPLE = 16'h6b2f;
		648: SAMPLE = 16'h6b4a;
		649: SAMPLE = 16'h6b66;
		650: SAMPLE = 16'h6b81;
		651: SAMPLE = 16'h6b9c;
		652: SAMPLE = 16'h6bb8;
		653: SAMPLE = 16'h6bd3;
		654: SAMPLE = 16'h6bee;
		655: SAMPLE = 16'h6c09;
		656: SAMPLE = 16'h6c24;
		657: SAMPLE = 16'h6c3f;
		658: SAMPLE = 16'h6c59;
		659: SAMPLE = 16'h6c74;
		660: SAMPLE = 16'h6c8f;
		661: SAMPLE = 16'h6ca9;
		662: SAMPLE = 16'h6cc4;
		663: SAMPLE = 16'h6cde;
		664: SAMPLE = 16'h6cf9;
		665: SAMPLE = 16'h6d13;
		666: SAMPLE = 16'h6d2d;
		667: SAMPLE = 16'h6d48;
		668: SAMPLE = 16'h6d62;
		669: SAMPLE = 16'h6d7c;
		670: SAMPLE = 16'h6d96;
		671: SAMPLE = 16'h6db0;
		672: SAMPLE = 16'h6dca;
		673: SAMPLE = 16'h6de3;
		674: SAMPLE = 16'h6dfd;
		675: SAMPLE = 16'h6e17;
		676: SAMPLE = 16'h6e30;
		677: SAMPLE = 16'h6e4a;
		678: SAMPLE = 16'h6e63;
		679: SAMPLE = 16'h6e7d;
		680: SAMPLE = 16'h6e96;
		681: SAMPLE = 16'h6eaf;
		682: SAMPLE = 16'h6ec9;
		683: SAMPLE = 16'h6ee2;
		684: SAMPLE = 16'h6efb;
		685: SAMPLE = 16'h6f14;
		686: SAMPLE = 16'h6f2d;
		687: SAMPLE = 16'h6f46;
		688: SAMPLE = 16'h6f5f;
		689: SAMPLE = 16'h6f77;
		690: SAMPLE = 16'h6f90;
		691: SAMPLE = 16'h6fa9;
		692: SAMPLE = 16'h6fc1;
		693: SAMPLE = 16'h6fda;
		694: SAMPLE = 16'h6ff2;
		695: SAMPLE = 16'h700a;
		696: SAMPLE = 16'h7023;
		697: SAMPLE = 16'h703b;
		698: SAMPLE = 16'h7053;
		699: SAMPLE = 16'h706b;
		700: SAMPLE = 16'h7083;
		701: SAMPLE = 16'h709b;
		702: SAMPLE = 16'h70b3;
		703: SAMPLE = 16'h70cb;
		704: SAMPLE = 16'h70e2;
		705: SAMPLE = 16'h70fa;
		706: SAMPLE = 16'h7112;
		707: SAMPLE = 16'h7129;
		708: SAMPLE = 16'h7141;
		709: SAMPLE = 16'h7158;
		710: SAMPLE = 16'h716f;
		711: SAMPLE = 16'h7186;
		712: SAMPLE = 16'h719e;
		713: SAMPLE = 16'h71b5;
		714: SAMPLE = 16'h71cc;
		715: SAMPLE = 16'h71e3;
		716: SAMPLE = 16'h71fa;
		717: SAMPLE = 16'h7211;
		718: SAMPLE = 16'h7227;
		719: SAMPLE = 16'h723e;
		720: SAMPLE = 16'h7255;
		721: SAMPLE = 16'h726b;
		722: SAMPLE = 16'h7282;
		723: SAMPLE = 16'h7298;
		724: SAMPLE = 16'h72af;
		725: SAMPLE = 16'h72c5;
		726: SAMPLE = 16'h72db;
		727: SAMPLE = 16'h72f1;
		728: SAMPLE = 16'h7307;
		729: SAMPLE = 16'h731d;
		730: SAMPLE = 16'h7333;
		731: SAMPLE = 16'h7349;
		732: SAMPLE = 16'h735f;
		733: SAMPLE = 16'h7375;
		734: SAMPLE = 16'h738a;
		735: SAMPLE = 16'h73a0;
		736: SAMPLE = 16'h73b5;
		737: SAMPLE = 16'h73cb;
		738: SAMPLE = 16'h73e0;
		739: SAMPLE = 16'h73f6;
		740: SAMPLE = 16'h740b;
		741: SAMPLE = 16'h7420;
		742: SAMPLE = 16'h7435;
		743: SAMPLE = 16'h744a;
		744: SAMPLE = 16'h745f;
		745: SAMPLE = 16'h7474;
		746: SAMPLE = 16'h7489;
		747: SAMPLE = 16'h749e;
		748: SAMPLE = 16'h74b2;
		749: SAMPLE = 16'h74c7;
		750: SAMPLE = 16'h74db;
		751: SAMPLE = 16'h74f0;
		752: SAMPLE = 16'h7504;
		753: SAMPLE = 16'h7519;
		754: SAMPLE = 16'h752d;
		755: SAMPLE = 16'h7541;
		756: SAMPLE = 16'h7555;
		757: SAMPLE = 16'h7569;
		758: SAMPLE = 16'h757d;
		759: SAMPLE = 16'h7591;
		760: SAMPLE = 16'h75a5;
		761: SAMPLE = 16'h75b9;
		762: SAMPLE = 16'h75cc;
		763: SAMPLE = 16'h75e0;
		764: SAMPLE = 16'h75f4;
		765: SAMPLE = 16'h7607;
		766: SAMPLE = 16'h761b;
		767: SAMPLE = 16'h762e;
		768: SAMPLE = 16'h7641;
		769: SAMPLE = 16'h7654;
		770: SAMPLE = 16'h7668;
		771: SAMPLE = 16'h767b;
		772: SAMPLE = 16'h768e;
		773: SAMPLE = 16'h76a0;
		774: SAMPLE = 16'h76b3;
		775: SAMPLE = 16'h76c6;
		776: SAMPLE = 16'h76d9;
		777: SAMPLE = 16'h76eb;
		778: SAMPLE = 16'h76fe;
		779: SAMPLE = 16'h7710;
		780: SAMPLE = 16'h7723;
		781: SAMPLE = 16'h7735;
		782: SAMPLE = 16'h7747;
		783: SAMPLE = 16'h775a;
		784: SAMPLE = 16'h776c;
		785: SAMPLE = 16'h777e;
		786: SAMPLE = 16'h7790;
		787: SAMPLE = 16'h77a2;
		788: SAMPLE = 16'h77b4;
		789: SAMPLE = 16'h77c5;
		790: SAMPLE = 16'h77d7;
		791: SAMPLE = 16'h77e9;
		792: SAMPLE = 16'h77fa;
		793: SAMPLE = 16'h780c;
		794: SAMPLE = 16'h781d;
		795: SAMPLE = 16'h782e;
		796: SAMPLE = 16'h7840;
		797: SAMPLE = 16'h7851;
		798: SAMPLE = 16'h7862;
		799: SAMPLE = 16'h7873;
		800: SAMPLE = 16'h7884;
		801: SAMPLE = 16'h7895;
		802: SAMPLE = 16'h78a6;
		803: SAMPLE = 16'h78b6;
		804: SAMPLE = 16'h78c7;
		805: SAMPLE = 16'h78d8;
		806: SAMPLE = 16'h78e8;
		807: SAMPLE = 16'h78f9;
		808: SAMPLE = 16'h7909;
		809: SAMPLE = 16'h7919;
		810: SAMPLE = 16'h792a;
		811: SAMPLE = 16'h793a;
		812: SAMPLE = 16'h794a;
		813: SAMPLE = 16'h795a;
		814: SAMPLE = 16'h796a;
		815: SAMPLE = 16'h797a;
		816: SAMPLE = 16'h798a;
		817: SAMPLE = 16'h7999;
		818: SAMPLE = 16'h79a9;
		819: SAMPLE = 16'h79b9;
		820: SAMPLE = 16'h79c8;
		821: SAMPLE = 16'h79d8;
		822: SAMPLE = 16'h79e7;
		823: SAMPLE = 16'h79f6;
		824: SAMPLE = 16'h7a05;
		825: SAMPLE = 16'h7a15;
		826: SAMPLE = 16'h7a24;
		827: SAMPLE = 16'h7a33;
		828: SAMPLE = 16'h7a42;
		829: SAMPLE = 16'h7a50;
		830: SAMPLE = 16'h7a5f;
		831: SAMPLE = 16'h7a6e;
		832: SAMPLE = 16'h7a7d;
		833: SAMPLE = 16'h7a8b;
		834: SAMPLE = 16'h7a9a;
		835: SAMPLE = 16'h7aa8;
		836: SAMPLE = 16'h7ab6;
		837: SAMPLE = 16'h7ac5;
		838: SAMPLE = 16'h7ad3;
		839: SAMPLE = 16'h7ae1;
		840: SAMPLE = 16'h7aef;
		841: SAMPLE = 16'h7afd;
		842: SAMPLE = 16'h7b0b;
		843: SAMPLE = 16'h7b19;
		844: SAMPLE = 16'h7b26;
		845: SAMPLE = 16'h7b34;
		846: SAMPLE = 16'h7b42;
		847: SAMPLE = 16'h7b4f;
		848: SAMPLE = 16'h7b5d;
		849: SAMPLE = 16'h7b6a;
		850: SAMPLE = 16'h7b77;
		851: SAMPLE = 16'h7b84;
		852: SAMPLE = 16'h7b92;
		853: SAMPLE = 16'h7b9f;
		854: SAMPLE = 16'h7bac;
		855: SAMPLE = 16'h7bb9;
		856: SAMPLE = 16'h7bc5;
		857: SAMPLE = 16'h7bd2;
		858: SAMPLE = 16'h7bdf;
		859: SAMPLE = 16'h7beb;
		860: SAMPLE = 16'h7bf8;
		861: SAMPLE = 16'h7c05;
		862: SAMPLE = 16'h7c11;
		863: SAMPLE = 16'h7c1d;
		864: SAMPLE = 16'h7c29;
		865: SAMPLE = 16'h7c36;
		866: SAMPLE = 16'h7c42;
		867: SAMPLE = 16'h7c4e;
		868: SAMPLE = 16'h7c5a;
		869: SAMPLE = 16'h7c66;
		870: SAMPLE = 16'h7c71;
		871: SAMPLE = 16'h7c7d;
		872: SAMPLE = 16'h7c89;
		873: SAMPLE = 16'h7c94;
		874: SAMPLE = 16'h7ca0;
		875: SAMPLE = 16'h7cab;
		876: SAMPLE = 16'h7cb7;
		877: SAMPLE = 16'h7cc2;
		878: SAMPLE = 16'h7ccd;
		879: SAMPLE = 16'h7cd8;
		880: SAMPLE = 16'h7ce3;
		881: SAMPLE = 16'h7cee;
		882: SAMPLE = 16'h7cf9;
		883: SAMPLE = 16'h7d04;
		884: SAMPLE = 16'h7d0f;
		885: SAMPLE = 16'h7d19;
		886: SAMPLE = 16'h7d24;
		887: SAMPLE = 16'h7d2f;
		888: SAMPLE = 16'h7d39;
		889: SAMPLE = 16'h7d43;
		890: SAMPLE = 16'h7d4e;
		891: SAMPLE = 16'h7d58;
		892: SAMPLE = 16'h7d62;
		893: SAMPLE = 16'h7d6c;
		894: SAMPLE = 16'h7d76;
		895: SAMPLE = 16'h7d80;
		896: SAMPLE = 16'h7d8a;
		897: SAMPLE = 16'h7d94;
		898: SAMPLE = 16'h7d9d;
		899: SAMPLE = 16'h7da7;
		900: SAMPLE = 16'h7db0;
		901: SAMPLE = 16'h7dba;
		902: SAMPLE = 16'h7dc3;
		903: SAMPLE = 16'h7dcd;
		904: SAMPLE = 16'h7dd6;
		905: SAMPLE = 16'h7ddf;
		906: SAMPLE = 16'h7de8;
		907: SAMPLE = 16'h7df1;
		908: SAMPLE = 16'h7dfa;
		909: SAMPLE = 16'h7e03;
		910: SAMPLE = 16'h7e0c;
		911: SAMPLE = 16'h7e14;
		912: SAMPLE = 16'h7e1d;
		913: SAMPLE = 16'h7e26;
		914: SAMPLE = 16'h7e2e;
		915: SAMPLE = 16'h7e37;
		916: SAMPLE = 16'h7e3f;
		917: SAMPLE = 16'h7e47;
		918: SAMPLE = 16'h7e4f;
		919: SAMPLE = 16'h7e57;
		920: SAMPLE = 16'h7e5f;
		921: SAMPLE = 16'h7e67;
		922: SAMPLE = 16'h7e6f;
		923: SAMPLE = 16'h7e77;
		924: SAMPLE = 16'h7e7f;
		925: SAMPLE = 16'h7e86;
		926: SAMPLE = 16'h7e8e;
		927: SAMPLE = 16'h7e95;
		928: SAMPLE = 16'h7e9d;
		929: SAMPLE = 16'h7ea4;
		930: SAMPLE = 16'h7eab;
		931: SAMPLE = 16'h7eb3;
		932: SAMPLE = 16'h7eba;
		933: SAMPLE = 16'h7ec1;
		934: SAMPLE = 16'h7ec8;
		935: SAMPLE = 16'h7ecf;
		936: SAMPLE = 16'h7ed5;
		937: SAMPLE = 16'h7edc;
		938: SAMPLE = 16'h7ee3;
		939: SAMPLE = 16'h7ee9;
		940: SAMPLE = 16'h7ef0;
		941: SAMPLE = 16'h7ef6;
		942: SAMPLE = 16'h7efd;
		943: SAMPLE = 16'h7f03;
		944: SAMPLE = 16'h7f09;
		945: SAMPLE = 16'h7f0f;
		946: SAMPLE = 16'h7f15;
		947: SAMPLE = 16'h7f1b;
		948: SAMPLE = 16'h7f21;
		949: SAMPLE = 16'h7f27;
		950: SAMPLE = 16'h7f2d;
		951: SAMPLE = 16'h7f32;
		952: SAMPLE = 16'h7f38;
		953: SAMPLE = 16'h7f3d;
		954: SAMPLE = 16'h7f43;
		955: SAMPLE = 16'h7f48;
		956: SAMPLE = 16'h7f4d;
		957: SAMPLE = 16'h7f53;
		958: SAMPLE = 16'h7f58;
		959: SAMPLE = 16'h7f5d;
		960: SAMPLE = 16'h7f62;
		961: SAMPLE = 16'h7f67;
		962: SAMPLE = 16'h7f6b;
		963: SAMPLE = 16'h7f70;
		964: SAMPLE = 16'h7f75;
		965: SAMPLE = 16'h7f79;
		966: SAMPLE = 16'h7f7e;
		967: SAMPLE = 16'h7f82;
		968: SAMPLE = 16'h7f87;
		969: SAMPLE = 16'h7f8b;
		970: SAMPLE = 16'h7f8f;
		971: SAMPLE = 16'h7f93;
		972: SAMPLE = 16'h7f97;
		973: SAMPLE = 16'h7f9b;
		974: SAMPLE = 16'h7f9f;
		975: SAMPLE = 16'h7fa3;
		976: SAMPLE = 16'h7fa7;
		977: SAMPLE = 16'h7faa;
		978: SAMPLE = 16'h7fae;
		979: SAMPLE = 16'h7fb1;
		980: SAMPLE = 16'h7fb5;
		981: SAMPLE = 16'h7fb8;
		982: SAMPLE = 16'h7fbc;
		983: SAMPLE = 16'h7fbf;
		984: SAMPLE = 16'h7fc2;
		985: SAMPLE = 16'h7fc5;
		986: SAMPLE = 16'h7fc8;
		987: SAMPLE = 16'h7fcb;
		988: SAMPLE = 16'h7fce;
		989: SAMPLE = 16'h7fd0;
		990: SAMPLE = 16'h7fd3;
		991: SAMPLE = 16'h7fd6;
		992: SAMPLE = 16'h7fd8;
		993: SAMPLE = 16'h7fda;
		994: SAMPLE = 16'h7fdd;
		995: SAMPLE = 16'h7fdf;
		996: SAMPLE = 16'h7fe1;
		997: SAMPLE = 16'h7fe3;
		998: SAMPLE = 16'h7fe5;
		999: SAMPLE = 16'h7fe7;
		1000: SAMPLE = 16'h7fe9;
		1001: SAMPLE = 16'h7feb;
		1002: SAMPLE = 16'h7fed;
		1003: SAMPLE = 16'h7fee;
		1004: SAMPLE = 16'h7ff0;
		1005: SAMPLE = 16'h7ff2;
		1006: SAMPLE = 16'h7ff3;
		1007: SAMPLE = 16'h7ff4;
		1008: SAMPLE = 16'h7ff6;
		1009: SAMPLE = 16'h7ff7;
		1010: SAMPLE = 16'h7ff8;
		1011: SAMPLE = 16'h7ff9;
		1012: SAMPLE = 16'h7ffa;
		1013: SAMPLE = 16'h7ffb;
		1014: SAMPLE = 16'h7ffc;
		1015: SAMPLE = 16'h7ffc;
		1016: SAMPLE = 16'h7ffd;
		1017: SAMPLE = 16'h7ffe;
		1018: SAMPLE = 16'h7ffe;
		1019: SAMPLE = 16'h7fff;
		1020: SAMPLE = 16'h7fff;
		1021: SAMPLE = 16'h7fff;
		1022: SAMPLE = 16'h7fff;
		1023: SAMPLE = 16'h7fff;
		1024: SAMPLE = 16'h8000;
		1025: SAMPLE = 16'h7fff;
		1026: SAMPLE = 16'h7fff;
		1027: SAMPLE = 16'h7fff;
		1028: SAMPLE = 16'h7fff;
		1029: SAMPLE = 16'h7fff;
		1030: SAMPLE = 16'h7ffe;
		1031: SAMPLE = 16'h7ffe;
		1032: SAMPLE = 16'h7ffd;
		1033: SAMPLE = 16'h7ffc;
		1034: SAMPLE = 16'h7ffc;
		1035: SAMPLE = 16'h7ffb;
		1036: SAMPLE = 16'h7ffa;
		1037: SAMPLE = 16'h7ff9;
		1038: SAMPLE = 16'h7ff8;
		1039: SAMPLE = 16'h7ff7;
		1040: SAMPLE = 16'h7ff6;
		1041: SAMPLE = 16'h7ff4;
		1042: SAMPLE = 16'h7ff3;
		1043: SAMPLE = 16'h7ff2;
		1044: SAMPLE = 16'h7ff0;
		1045: SAMPLE = 16'h7fee;
		1046: SAMPLE = 16'h7fed;
		1047: SAMPLE = 16'h7feb;
		1048: SAMPLE = 16'h7fe9;
		1049: SAMPLE = 16'h7fe7;
		1050: SAMPLE = 16'h7fe5;
		1051: SAMPLE = 16'h7fe3;
		1052: SAMPLE = 16'h7fe1;
		1053: SAMPLE = 16'h7fdf;
		1054: SAMPLE = 16'h7fdd;
		1055: SAMPLE = 16'h7fda;
		1056: SAMPLE = 16'h7fd8;
		1057: SAMPLE = 16'h7fd6;
		1058: SAMPLE = 16'h7fd3;
		1059: SAMPLE = 16'h7fd0;
		1060: SAMPLE = 16'h7fce;
		1061: SAMPLE = 16'h7fcb;
		1062: SAMPLE = 16'h7fc8;
		1063: SAMPLE = 16'h7fc5;
		1064: SAMPLE = 16'h7fc2;
		1065: SAMPLE = 16'h7fbf;
		1066: SAMPLE = 16'h7fbc;
		1067: SAMPLE = 16'h7fb8;
		1068: SAMPLE = 16'h7fb5;
		1069: SAMPLE = 16'h7fb1;
		1070: SAMPLE = 16'h7fae;
		1071: SAMPLE = 16'h7faa;
		1072: SAMPLE = 16'h7fa7;
		1073: SAMPLE = 16'h7fa3;
		1074: SAMPLE = 16'h7f9f;
		1075: SAMPLE = 16'h7f9b;
		1076: SAMPLE = 16'h7f97;
		1077: SAMPLE = 16'h7f93;
		1078: SAMPLE = 16'h7f8f;
		1079: SAMPLE = 16'h7f8b;
		1080: SAMPLE = 16'h7f87;
		1081: SAMPLE = 16'h7f82;
		1082: SAMPLE = 16'h7f7e;
		1083: SAMPLE = 16'h7f79;
		1084: SAMPLE = 16'h7f75;
		1085: SAMPLE = 16'h7f70;
		1086: SAMPLE = 16'h7f6b;
		1087: SAMPLE = 16'h7f67;
		1088: SAMPLE = 16'h7f62;
		1089: SAMPLE = 16'h7f5d;
		1090: SAMPLE = 16'h7f58;
		1091: SAMPLE = 16'h7f53;
		1092: SAMPLE = 16'h7f4d;
		1093: SAMPLE = 16'h7f48;
		1094: SAMPLE = 16'h7f43;
		1095: SAMPLE = 16'h7f3d;
		1096: SAMPLE = 16'h7f38;
		1097: SAMPLE = 16'h7f32;
		1098: SAMPLE = 16'h7f2d;
		1099: SAMPLE = 16'h7f27;
		1100: SAMPLE = 16'h7f21;
		1101: SAMPLE = 16'h7f1b;
		1102: SAMPLE = 16'h7f15;
		1103: SAMPLE = 16'h7f0f;
		1104: SAMPLE = 16'h7f09;
		1105: SAMPLE = 16'h7f03;
		1106: SAMPLE = 16'h7efd;
		1107: SAMPLE = 16'h7ef6;
		1108: SAMPLE = 16'h7ef0;
		1109: SAMPLE = 16'h7ee9;
		1110: SAMPLE = 16'h7ee3;
		1111: SAMPLE = 16'h7edc;
		1112: SAMPLE = 16'h7ed5;
		1113: SAMPLE = 16'h7ecf;
		1114: SAMPLE = 16'h7ec8;
		1115: SAMPLE = 16'h7ec1;
		1116: SAMPLE = 16'h7eba;
		1117: SAMPLE = 16'h7eb3;
		1118: SAMPLE = 16'h7eab;
		1119: SAMPLE = 16'h7ea4;
		1120: SAMPLE = 16'h7e9d;
		1121: SAMPLE = 16'h7e95;
		1122: SAMPLE = 16'h7e8e;
		1123: SAMPLE = 16'h7e86;
		1124: SAMPLE = 16'h7e7f;
		1125: SAMPLE = 16'h7e77;
		1126: SAMPLE = 16'h7e6f;
		1127: SAMPLE = 16'h7e67;
		1128: SAMPLE = 16'h7e5f;
		1129: SAMPLE = 16'h7e57;
		1130: SAMPLE = 16'h7e4f;
		1131: SAMPLE = 16'h7e47;
		1132: SAMPLE = 16'h7e3f;
		1133: SAMPLE = 16'h7e37;
		1134: SAMPLE = 16'h7e2e;
		1135: SAMPLE = 16'h7e26;
		1136: SAMPLE = 16'h7e1d;
		1137: SAMPLE = 16'h7e14;
		1138: SAMPLE = 16'h7e0c;
		1139: SAMPLE = 16'h7e03;
		1140: SAMPLE = 16'h7dfa;
		1141: SAMPLE = 16'h7df1;
		1142: SAMPLE = 16'h7de8;
		1143: SAMPLE = 16'h7ddf;
		1144: SAMPLE = 16'h7dd6;
		1145: SAMPLE = 16'h7dcd;
		1146: SAMPLE = 16'h7dc3;
		1147: SAMPLE = 16'h7dba;
		1148: SAMPLE = 16'h7db0;
		1149: SAMPLE = 16'h7da7;
		1150: SAMPLE = 16'h7d9d;
		1151: SAMPLE = 16'h7d94;
		1152: SAMPLE = 16'h7d8a;
		1153: SAMPLE = 16'h7d80;
		1154: SAMPLE = 16'h7d76;
		1155: SAMPLE = 16'h7d6c;
		1156: SAMPLE = 16'h7d62;
		1157: SAMPLE = 16'h7d58;
		1158: SAMPLE = 16'h7d4e;
		1159: SAMPLE = 16'h7d43;
		1160: SAMPLE = 16'h7d39;
		1161: SAMPLE = 16'h7d2f;
		1162: SAMPLE = 16'h7d24;
		1163: SAMPLE = 16'h7d19;
		1164: SAMPLE = 16'h7d0f;
		1165: SAMPLE = 16'h7d04;
		1166: SAMPLE = 16'h7cf9;
		1167: SAMPLE = 16'h7cee;
		1168: SAMPLE = 16'h7ce3;
		1169: SAMPLE = 16'h7cd8;
		1170: SAMPLE = 16'h7ccd;
		1171: SAMPLE = 16'h7cc2;
		1172: SAMPLE = 16'h7cb7;
		1173: SAMPLE = 16'h7cab;
		1174: SAMPLE = 16'h7ca0;
		1175: SAMPLE = 16'h7c94;
		1176: SAMPLE = 16'h7c89;
		1177: SAMPLE = 16'h7c7d;
		1178: SAMPLE = 16'h7c71;
		1179: SAMPLE = 16'h7c66;
		1180: SAMPLE = 16'h7c5a;
		1181: SAMPLE = 16'h7c4e;
		1182: SAMPLE = 16'h7c42;
		1183: SAMPLE = 16'h7c36;
		1184: SAMPLE = 16'h7c29;
		1185: SAMPLE = 16'h7c1d;
		1186: SAMPLE = 16'h7c11;
		1187: SAMPLE = 16'h7c05;
		1188: SAMPLE = 16'h7bf8;
		1189: SAMPLE = 16'h7beb;
		1190: SAMPLE = 16'h7bdf;
		1191: SAMPLE = 16'h7bd2;
		1192: SAMPLE = 16'h7bc5;
		1193: SAMPLE = 16'h7bb9;
		1194: SAMPLE = 16'h7bac;
		1195: SAMPLE = 16'h7b9f;
		1196: SAMPLE = 16'h7b92;
		1197: SAMPLE = 16'h7b84;
		1198: SAMPLE = 16'h7b77;
		1199: SAMPLE = 16'h7b6a;
		1200: SAMPLE = 16'h7b5d;
		1201: SAMPLE = 16'h7b4f;
		1202: SAMPLE = 16'h7b42;
		1203: SAMPLE = 16'h7b34;
		1204: SAMPLE = 16'h7b26;
		1205: SAMPLE = 16'h7b19;
		1206: SAMPLE = 16'h7b0b;
		1207: SAMPLE = 16'h7afd;
		1208: SAMPLE = 16'h7aef;
		1209: SAMPLE = 16'h7ae1;
		1210: SAMPLE = 16'h7ad3;
		1211: SAMPLE = 16'h7ac5;
		1212: SAMPLE = 16'h7ab6;
		1213: SAMPLE = 16'h7aa8;
		1214: SAMPLE = 16'h7a9a;
		1215: SAMPLE = 16'h7a8b;
		1216: SAMPLE = 16'h7a7d;
		1217: SAMPLE = 16'h7a6e;
		1218: SAMPLE = 16'h7a5f;
		1219: SAMPLE = 16'h7a50;
		1220: SAMPLE = 16'h7a42;
		1221: SAMPLE = 16'h7a33;
		1222: SAMPLE = 16'h7a24;
		1223: SAMPLE = 16'h7a15;
		1224: SAMPLE = 16'h7a05;
		1225: SAMPLE = 16'h79f6;
		1226: SAMPLE = 16'h79e7;
		1227: SAMPLE = 16'h79d8;
		1228: SAMPLE = 16'h79c8;
		1229: SAMPLE = 16'h79b9;
		1230: SAMPLE = 16'h79a9;
		1231: SAMPLE = 16'h7999;
		1232: SAMPLE = 16'h798a;
		1233: SAMPLE = 16'h797a;
		1234: SAMPLE = 16'h796a;
		1235: SAMPLE = 16'h795a;
		1236: SAMPLE = 16'h794a;
		1237: SAMPLE = 16'h793a;
		1238: SAMPLE = 16'h792a;
		1239: SAMPLE = 16'h7919;
		1240: SAMPLE = 16'h7909;
		1241: SAMPLE = 16'h78f9;
		1242: SAMPLE = 16'h78e8;
		1243: SAMPLE = 16'h78d8;
		1244: SAMPLE = 16'h78c7;
		1245: SAMPLE = 16'h78b6;
		1246: SAMPLE = 16'h78a6;
		1247: SAMPLE = 16'h7895;
		1248: SAMPLE = 16'h7884;
		1249: SAMPLE = 16'h7873;
		1250: SAMPLE = 16'h7862;
		1251: SAMPLE = 16'h7851;
		1252: SAMPLE = 16'h7840;
		1253: SAMPLE = 16'h782e;
		1254: SAMPLE = 16'h781d;
		1255: SAMPLE = 16'h780c;
		1256: SAMPLE = 16'h77fa;
		1257: SAMPLE = 16'h77e9;
		1258: SAMPLE = 16'h77d7;
		1259: SAMPLE = 16'h77c5;
		1260: SAMPLE = 16'h77b4;
		1261: SAMPLE = 16'h77a2;
		1262: SAMPLE = 16'h7790;
		1263: SAMPLE = 16'h777e;
		1264: SAMPLE = 16'h776c;
		1265: SAMPLE = 16'h775a;
		1266: SAMPLE = 16'h7747;
		1267: SAMPLE = 16'h7735;
		1268: SAMPLE = 16'h7723;
		1269: SAMPLE = 16'h7710;
		1270: SAMPLE = 16'h76fe;
		1271: SAMPLE = 16'h76eb;
		1272: SAMPLE = 16'h76d9;
		1273: SAMPLE = 16'h76c6;
		1274: SAMPLE = 16'h76b3;
		1275: SAMPLE = 16'h76a0;
		1276: SAMPLE = 16'h768e;
		1277: SAMPLE = 16'h767b;
		1278: SAMPLE = 16'h7668;
		1279: SAMPLE = 16'h7654;
		1280: SAMPLE = 16'h7641;
		1281: SAMPLE = 16'h762e;
		1282: SAMPLE = 16'h761b;
		1283: SAMPLE = 16'h7607;
		1284: SAMPLE = 16'h75f4;
		1285: SAMPLE = 16'h75e0;
		1286: SAMPLE = 16'h75cc;
		1287: SAMPLE = 16'h75b9;
		1288: SAMPLE = 16'h75a5;
		1289: SAMPLE = 16'h7591;
		1290: SAMPLE = 16'h757d;
		1291: SAMPLE = 16'h7569;
		1292: SAMPLE = 16'h7555;
		1293: SAMPLE = 16'h7541;
		1294: SAMPLE = 16'h752d;
		1295: SAMPLE = 16'h7519;
		1296: SAMPLE = 16'h7504;
		1297: SAMPLE = 16'h74f0;
		1298: SAMPLE = 16'h74db;
		1299: SAMPLE = 16'h74c7;
		1300: SAMPLE = 16'h74b2;
		1301: SAMPLE = 16'h749e;
		1302: SAMPLE = 16'h7489;
		1303: SAMPLE = 16'h7474;
		1304: SAMPLE = 16'h745f;
		1305: SAMPLE = 16'h744a;
		1306: SAMPLE = 16'h7435;
		1307: SAMPLE = 16'h7420;
		1308: SAMPLE = 16'h740b;
		1309: SAMPLE = 16'h73f6;
		1310: SAMPLE = 16'h73e0;
		1311: SAMPLE = 16'h73cb;
		1312: SAMPLE = 16'h73b5;
		1313: SAMPLE = 16'h73a0;
		1314: SAMPLE = 16'h738a;
		1315: SAMPLE = 16'h7375;
		1316: SAMPLE = 16'h735f;
		1317: SAMPLE = 16'h7349;
		1318: SAMPLE = 16'h7333;
		1319: SAMPLE = 16'h731d;
		1320: SAMPLE = 16'h7307;
		1321: SAMPLE = 16'h72f1;
		1322: SAMPLE = 16'h72db;
		1323: SAMPLE = 16'h72c5;
		1324: SAMPLE = 16'h72af;
		1325: SAMPLE = 16'h7298;
		1326: SAMPLE = 16'h7282;
		1327: SAMPLE = 16'h726b;
		1328: SAMPLE = 16'h7255;
		1329: SAMPLE = 16'h723e;
		1330: SAMPLE = 16'h7227;
		1331: SAMPLE = 16'h7211;
		1332: SAMPLE = 16'h71fa;
		1333: SAMPLE = 16'h71e3;
		1334: SAMPLE = 16'h71cc;
		1335: SAMPLE = 16'h71b5;
		1336: SAMPLE = 16'h719e;
		1337: SAMPLE = 16'h7186;
		1338: SAMPLE = 16'h716f;
		1339: SAMPLE = 16'h7158;
		1340: SAMPLE = 16'h7141;
		1341: SAMPLE = 16'h7129;
		1342: SAMPLE = 16'h7112;
		1343: SAMPLE = 16'h70fa;
		1344: SAMPLE = 16'h70e2;
		1345: SAMPLE = 16'h70cb;
		1346: SAMPLE = 16'h70b3;
		1347: SAMPLE = 16'h709b;
		1348: SAMPLE = 16'h7083;
		1349: SAMPLE = 16'h706b;
		1350: SAMPLE = 16'h7053;
		1351: SAMPLE = 16'h703b;
		1352: SAMPLE = 16'h7023;
		1353: SAMPLE = 16'h700a;
		1354: SAMPLE = 16'h6ff2;
		1355: SAMPLE = 16'h6fda;
		1356: SAMPLE = 16'h6fc1;
		1357: SAMPLE = 16'h6fa9;
		1358: SAMPLE = 16'h6f90;
		1359: SAMPLE = 16'h6f77;
		1360: SAMPLE = 16'h6f5f;
		1361: SAMPLE = 16'h6f46;
		1362: SAMPLE = 16'h6f2d;
		1363: SAMPLE = 16'h6f14;
		1364: SAMPLE = 16'h6efb;
		1365: SAMPLE = 16'h6ee2;
		1366: SAMPLE = 16'h6ec9;
		1367: SAMPLE = 16'h6eaf;
		1368: SAMPLE = 16'h6e96;
		1369: SAMPLE = 16'h6e7d;
		1370: SAMPLE = 16'h6e63;
		1371: SAMPLE = 16'h6e4a;
		1372: SAMPLE = 16'h6e30;
		1373: SAMPLE = 16'h6e17;
		1374: SAMPLE = 16'h6dfd;
		1375: SAMPLE = 16'h6de3;
		1376: SAMPLE = 16'h6dca;
		1377: SAMPLE = 16'h6db0;
		1378: SAMPLE = 16'h6d96;
		1379: SAMPLE = 16'h6d7c;
		1380: SAMPLE = 16'h6d62;
		1381: SAMPLE = 16'h6d48;
		1382: SAMPLE = 16'h6d2d;
		1383: SAMPLE = 16'h6d13;
		1384: SAMPLE = 16'h6cf9;
		1385: SAMPLE = 16'h6cde;
		1386: SAMPLE = 16'h6cc4;
		1387: SAMPLE = 16'h6ca9;
		1388: SAMPLE = 16'h6c8f;
		1389: SAMPLE = 16'h6c74;
		1390: SAMPLE = 16'h6c59;
		1391: SAMPLE = 16'h6c3f;
		1392: SAMPLE = 16'h6c24;
		1393: SAMPLE = 16'h6c09;
		1394: SAMPLE = 16'h6bee;
		1395: SAMPLE = 16'h6bd3;
		1396: SAMPLE = 16'h6bb8;
		1397: SAMPLE = 16'h6b9c;
		1398: SAMPLE = 16'h6b81;
		1399: SAMPLE = 16'h6b66;
		1400: SAMPLE = 16'h6b4a;
		1401: SAMPLE = 16'h6b2f;
		1402: SAMPLE = 16'h6b13;
		1403: SAMPLE = 16'h6af8;
		1404: SAMPLE = 16'h6adc;
		1405: SAMPLE = 16'h6ac1;
		1406: SAMPLE = 16'h6aa5;
		1407: SAMPLE = 16'h6a89;
		1408: SAMPLE = 16'h6a6d;
		1409: SAMPLE = 16'h6a51;
		1410: SAMPLE = 16'h6a35;
		1411: SAMPLE = 16'h6a19;
		1412: SAMPLE = 16'h69fd;
		1413: SAMPLE = 16'h69e1;
		1414: SAMPLE = 16'h69c4;
		1415: SAMPLE = 16'h69a8;
		1416: SAMPLE = 16'h698c;
		1417: SAMPLE = 16'h696f;
		1418: SAMPLE = 16'h6953;
		1419: SAMPLE = 16'h6936;
		1420: SAMPLE = 16'h6919;
		1421: SAMPLE = 16'h68fd;
		1422: SAMPLE = 16'h68e0;
		1423: SAMPLE = 16'h68c3;
		1424: SAMPLE = 16'h68a6;
		1425: SAMPLE = 16'h6889;
		1426: SAMPLE = 16'h686c;
		1427: SAMPLE = 16'h684f;
		1428: SAMPLE = 16'h6832;
		1429: SAMPLE = 16'h6815;
		1430: SAMPLE = 16'h67f7;
		1431: SAMPLE = 16'h67da;
		1432: SAMPLE = 16'h67bd;
		1433: SAMPLE = 16'h679f;
		1434: SAMPLE = 16'h6782;
		1435: SAMPLE = 16'h6764;
		1436: SAMPLE = 16'h6746;
		1437: SAMPLE = 16'h6729;
		1438: SAMPLE = 16'h670b;
		1439: SAMPLE = 16'h66ed;
		1440: SAMPLE = 16'h66cf;
		1441: SAMPLE = 16'h66b1;
		1442: SAMPLE = 16'h6693;
		1443: SAMPLE = 16'h6675;
		1444: SAMPLE = 16'h6657;
		1445: SAMPLE = 16'h6639;
		1446: SAMPLE = 16'h661a;
		1447: SAMPLE = 16'h65fc;
		1448: SAMPLE = 16'h65dd;
		1449: SAMPLE = 16'h65bf;
		1450: SAMPLE = 16'h65a0;
		1451: SAMPLE = 16'h6582;
		1452: SAMPLE = 16'h6563;
		1453: SAMPLE = 16'h6545;
		1454: SAMPLE = 16'h6526;
		1455: SAMPLE = 16'h6507;
		1456: SAMPLE = 16'h64e8;
		1457: SAMPLE = 16'h64c9;
		1458: SAMPLE = 16'h64aa;
		1459: SAMPLE = 16'h648b;
		1460: SAMPLE = 16'h646c;
		1461: SAMPLE = 16'h644d;
		1462: SAMPLE = 16'h642d;
		1463: SAMPLE = 16'h640e;
		1464: SAMPLE = 16'h63ef;
		1465: SAMPLE = 16'h63cf;
		1466: SAMPLE = 16'h63b0;
		1467: SAMPLE = 16'h6390;
		1468: SAMPLE = 16'h6371;
		1469: SAMPLE = 16'h6351;
		1470: SAMPLE = 16'h6331;
		1471: SAMPLE = 16'h6311;
		1472: SAMPLE = 16'h62f2;
		1473: SAMPLE = 16'h62d2;
		1474: SAMPLE = 16'h62b2;
		1475: SAMPLE = 16'h6292;
		1476: SAMPLE = 16'h6271;
		1477: SAMPLE = 16'h6251;
		1478: SAMPLE = 16'h6231;
		1479: SAMPLE = 16'h6211;
		1480: SAMPLE = 16'h61f1;
		1481: SAMPLE = 16'h61d0;
		1482: SAMPLE = 16'h61b0;
		1483: SAMPLE = 16'h618f;
		1484: SAMPLE = 16'h616f;
		1485: SAMPLE = 16'h614e;
		1486: SAMPLE = 16'h612d;
		1487: SAMPLE = 16'h610d;
		1488: SAMPLE = 16'h60ec;
		1489: SAMPLE = 16'h60cb;
		1490: SAMPLE = 16'h60aa;
		1491: SAMPLE = 16'h6089;
		1492: SAMPLE = 16'h6068;
		1493: SAMPLE = 16'h6047;
		1494: SAMPLE = 16'h6026;
		1495: SAMPLE = 16'h6004;
		1496: SAMPLE = 16'h5fe3;
		1497: SAMPLE = 16'h5fc2;
		1498: SAMPLE = 16'h5fa0;
		1499: SAMPLE = 16'h5f7f;
		1500: SAMPLE = 16'h5f5e;
		1501: SAMPLE = 16'h5f3c;
		1502: SAMPLE = 16'h5f1a;
		1503: SAMPLE = 16'h5ef9;
		1504: SAMPLE = 16'h5ed7;
		1505: SAMPLE = 16'h5eb5;
		1506: SAMPLE = 16'h5e93;
		1507: SAMPLE = 16'h5e71;
		1508: SAMPLE = 16'h5e50;
		1509: SAMPLE = 16'h5e2d;
		1510: SAMPLE = 16'h5e0b;
		1511: SAMPLE = 16'h5de9;
		1512: SAMPLE = 16'h5dc7;
		1513: SAMPLE = 16'h5da5;
		1514: SAMPLE = 16'h5d83;
		1515: SAMPLE = 16'h5d60;
		1516: SAMPLE = 16'h5d3e;
		1517: SAMPLE = 16'h5d1b;
		1518: SAMPLE = 16'h5cf9;
		1519: SAMPLE = 16'h5cd6;
		1520: SAMPLE = 16'h5cb4;
		1521: SAMPLE = 16'h5c91;
		1522: SAMPLE = 16'h5c6e;
		1523: SAMPLE = 16'h5c4b;
		1524: SAMPLE = 16'h5c29;
		1525: SAMPLE = 16'h5c06;
		1526: SAMPLE = 16'h5be3;
		1527: SAMPLE = 16'h5bc0;
		1528: SAMPLE = 16'h5b9d;
		1529: SAMPLE = 16'h5b79;
		1530: SAMPLE = 16'h5b56;
		1531: SAMPLE = 16'h5b33;
		1532: SAMPLE = 16'h5b10;
		1533: SAMPLE = 16'h5aec;
		1534: SAMPLE = 16'h5ac9;
		1535: SAMPLE = 16'h5aa5;
		1536: SAMPLE = 16'h5a82;
		1537: SAMPLE = 16'h5a5e;
		1538: SAMPLE = 16'h5a3b;
		1539: SAMPLE = 16'h5a17;
		1540: SAMPLE = 16'h59f3;
		1541: SAMPLE = 16'h59d0;
		1542: SAMPLE = 16'h59ac;
		1543: SAMPLE = 16'h5988;
		1544: SAMPLE = 16'h5964;
		1545: SAMPLE = 16'h5940;
		1546: SAMPLE = 16'h591c;
		1547: SAMPLE = 16'h58f8;
		1548: SAMPLE = 16'h58d4;
		1549: SAMPLE = 16'h58af;
		1550: SAMPLE = 16'h588b;
		1551: SAMPLE = 16'h5867;
		1552: SAMPLE = 16'h5842;
		1553: SAMPLE = 16'h581e;
		1554: SAMPLE = 16'h57f9;
		1555: SAMPLE = 16'h57d5;
		1556: SAMPLE = 16'h57b0;
		1557: SAMPLE = 16'h578c;
		1558: SAMPLE = 16'h5767;
		1559: SAMPLE = 16'h5742;
		1560: SAMPLE = 16'h571d;
		1561: SAMPLE = 16'h56f9;
		1562: SAMPLE = 16'h56d4;
		1563: SAMPLE = 16'h56af;
		1564: SAMPLE = 16'h568a;
		1565: SAMPLE = 16'h5665;
		1566: SAMPLE = 16'h5640;
		1567: SAMPLE = 16'h561a;
		1568: SAMPLE = 16'h55f5;
		1569: SAMPLE = 16'h55d0;
		1570: SAMPLE = 16'h55ab;
		1571: SAMPLE = 16'h5585;
		1572: SAMPLE = 16'h5560;
		1573: SAMPLE = 16'h553a;
		1574: SAMPLE = 16'h5515;
		1575: SAMPLE = 16'h54ef;
		1576: SAMPLE = 16'h54ca;
		1577: SAMPLE = 16'h54a4;
		1578: SAMPLE = 16'h547e;
		1579: SAMPLE = 16'h5458;
		1580: SAMPLE = 16'h5433;
		1581: SAMPLE = 16'h540d;
		1582: SAMPLE = 16'h53e7;
		1583: SAMPLE = 16'h53c1;
		1584: SAMPLE = 16'h539b;
		1585: SAMPLE = 16'h5375;
		1586: SAMPLE = 16'h534e;
		1587: SAMPLE = 16'h5328;
		1588: SAMPLE = 16'h5302;
		1589: SAMPLE = 16'h52dc;
		1590: SAMPLE = 16'h52b5;
		1591: SAMPLE = 16'h528f;
		1592: SAMPLE = 16'h5269;
		1593: SAMPLE = 16'h5242;
		1594: SAMPLE = 16'h521c;
		1595: SAMPLE = 16'h51f5;
		1596: SAMPLE = 16'h51ce;
		1597: SAMPLE = 16'h51a8;
		1598: SAMPLE = 16'h5181;
		1599: SAMPLE = 16'h515a;
		1600: SAMPLE = 16'h5133;
		1601: SAMPLE = 16'h510c;
		1602: SAMPLE = 16'h50e5;
		1603: SAMPLE = 16'h50bf;
		1604: SAMPLE = 16'h5097;
		1605: SAMPLE = 16'h5070;
		1606: SAMPLE = 16'h5049;
		1607: SAMPLE = 16'h5022;
		1608: SAMPLE = 16'h4ffb;
		1609: SAMPLE = 16'h4fd4;
		1610: SAMPLE = 16'h4fac;
		1611: SAMPLE = 16'h4f85;
		1612: SAMPLE = 16'h4f5e;
		1613: SAMPLE = 16'h4f36;
		1614: SAMPLE = 16'h4f0f;
		1615: SAMPLE = 16'h4ee7;
		1616: SAMPLE = 16'h4ebf;
		1617: SAMPLE = 16'h4e98;
		1618: SAMPLE = 16'h4e70;
		1619: SAMPLE = 16'h4e48;
		1620: SAMPLE = 16'h4e21;
		1621: SAMPLE = 16'h4df9;
		1622: SAMPLE = 16'h4dd1;
		1623: SAMPLE = 16'h4da9;
		1624: SAMPLE = 16'h4d81;
		1625: SAMPLE = 16'h4d59;
		1626: SAMPLE = 16'h4d31;
		1627: SAMPLE = 16'h4d09;
		1628: SAMPLE = 16'h4ce1;
		1629: SAMPLE = 16'h4cb8;
		1630: SAMPLE = 16'h4c90;
		1631: SAMPLE = 16'h4c68;
		1632: SAMPLE = 16'h4c3f;
		1633: SAMPLE = 16'h4c17;
		1634: SAMPLE = 16'h4bef;
		1635: SAMPLE = 16'h4bc6;
		1636: SAMPLE = 16'h4b9e;
		1637: SAMPLE = 16'h4b75;
		1638: SAMPLE = 16'h4b4c;
		1639: SAMPLE = 16'h4b24;
		1640: SAMPLE = 16'h4afb;
		1641: SAMPLE = 16'h4ad2;
		1642: SAMPLE = 16'h4aa9;
		1643: SAMPLE = 16'h4a81;
		1644: SAMPLE = 16'h4a58;
		1645: SAMPLE = 16'h4a2f;
		1646: SAMPLE = 16'h4a06;
		1647: SAMPLE = 16'h49dd;
		1648: SAMPLE = 16'h49b4;
		1649: SAMPLE = 16'h498a;
		1650: SAMPLE = 16'h4961;
		1651: SAMPLE = 16'h4938;
		1652: SAMPLE = 16'h490f;
		1653: SAMPLE = 16'h48e6;
		1654: SAMPLE = 16'h48bc;
		1655: SAMPLE = 16'h4893;
		1656: SAMPLE = 16'h4869;
		1657: SAMPLE = 16'h4840;
		1658: SAMPLE = 16'h4816;
		1659: SAMPLE = 16'h47ed;
		1660: SAMPLE = 16'h47c3;
		1661: SAMPLE = 16'h479a;
		1662: SAMPLE = 16'h4770;
		1663: SAMPLE = 16'h4746;
		1664: SAMPLE = 16'h471c;
		1665: SAMPLE = 16'h46f3;
		1666: SAMPLE = 16'h46c9;
		1667: SAMPLE = 16'h469f;
		1668: SAMPLE = 16'h4675;
		1669: SAMPLE = 16'h464b;
		1670: SAMPLE = 16'h4621;
		1671: SAMPLE = 16'h45f7;
		1672: SAMPLE = 16'h45cd;
		1673: SAMPLE = 16'h45a3;
		1674: SAMPLE = 16'h4578;
		1675: SAMPLE = 16'h454e;
		1676: SAMPLE = 16'h4524;
		1677: SAMPLE = 16'h44fa;
		1678: SAMPLE = 16'h44cf;
		1679: SAMPLE = 16'h44a5;
		1680: SAMPLE = 16'h447a;
		1681: SAMPLE = 16'h4450;
		1682: SAMPLE = 16'h4425;
		1683: SAMPLE = 16'h43fb;
		1684: SAMPLE = 16'h43d0;
		1685: SAMPLE = 16'h43a5;
		1686: SAMPLE = 16'h437b;
		1687: SAMPLE = 16'h4350;
		1688: SAMPLE = 16'h4325;
		1689: SAMPLE = 16'h42fa;
		1690: SAMPLE = 16'h42d0;
		1691: SAMPLE = 16'h42a5;
		1692: SAMPLE = 16'h427a;
		1693: SAMPLE = 16'h424f;
		1694: SAMPLE = 16'h4224;
		1695: SAMPLE = 16'h41f9;
		1696: SAMPLE = 16'h41ce;
		1697: SAMPLE = 16'h41a2;
		1698: SAMPLE = 16'h4177;
		1699: SAMPLE = 16'h414c;
		1700: SAMPLE = 16'h4121;
		1701: SAMPLE = 16'h40f6;
		1702: SAMPLE = 16'h40ca;
		1703: SAMPLE = 16'h409f;
		1704: SAMPLE = 16'h4073;
		1705: SAMPLE = 16'h4048;
		1706: SAMPLE = 16'h401d;
		1707: SAMPLE = 16'h3ff1;
		1708: SAMPLE = 16'h3fc5;
		1709: SAMPLE = 16'h3f9a;
		1710: SAMPLE = 16'h3f6e;
		1711: SAMPLE = 16'h3f43;
		1712: SAMPLE = 16'h3f17;
		1713: SAMPLE = 16'h3eeb;
		1714: SAMPLE = 16'h3ebf;
		1715: SAMPLE = 16'h3e93;
		1716: SAMPLE = 16'h3e68;
		1717: SAMPLE = 16'h3e3c;
		1718: SAMPLE = 16'h3e10;
		1719: SAMPLE = 16'h3de4;
		1720: SAMPLE = 16'h3db8;
		1721: SAMPLE = 16'h3d8c;
		1722: SAMPLE = 16'h3d60;
		1723: SAMPLE = 16'h3d33;
		1724: SAMPLE = 16'h3d07;
		1725: SAMPLE = 16'h3cdb;
		1726: SAMPLE = 16'h3caf;
		1727: SAMPLE = 16'h3c83;
		1728: SAMPLE = 16'h3c56;
		1729: SAMPLE = 16'h3c2a;
		1730: SAMPLE = 16'h3bfd;
		1731: SAMPLE = 16'h3bd1;
		1732: SAMPLE = 16'h3ba5;
		1733: SAMPLE = 16'h3b78;
		1734: SAMPLE = 16'h3b4c;
		1735: SAMPLE = 16'h3b1f;
		1736: SAMPLE = 16'h3af2;
		1737: SAMPLE = 16'h3ac6;
		1738: SAMPLE = 16'h3a99;
		1739: SAMPLE = 16'h3a6c;
		1740: SAMPLE = 16'h3a40;
		1741: SAMPLE = 16'h3a13;
		1742: SAMPLE = 16'h39e6;
		1743: SAMPLE = 16'h39b9;
		1744: SAMPLE = 16'h398c;
		1745: SAMPLE = 16'h395f;
		1746: SAMPLE = 16'h3932;
		1747: SAMPLE = 16'h3906;
		1748: SAMPLE = 16'h38d8;
		1749: SAMPLE = 16'h38ab;
		1750: SAMPLE = 16'h387e;
		1751: SAMPLE = 16'h3851;
		1752: SAMPLE = 16'h3824;
		1753: SAMPLE = 16'h37f7;
		1754: SAMPLE = 16'h37ca;
		1755: SAMPLE = 16'h379c;
		1756: SAMPLE = 16'h376f;
		1757: SAMPLE = 16'h3742;
		1758: SAMPLE = 16'h3714;
		1759: SAMPLE = 16'h36e7;
		1760: SAMPLE = 16'h36ba;
		1761: SAMPLE = 16'h368c;
		1762: SAMPLE = 16'h365f;
		1763: SAMPLE = 16'h3631;
		1764: SAMPLE = 16'h3604;
		1765: SAMPLE = 16'h35d6;
		1766: SAMPLE = 16'h35a8;
		1767: SAMPLE = 16'h357b;
		1768: SAMPLE = 16'h354d;
		1769: SAMPLE = 16'h351f;
		1770: SAMPLE = 16'h34f2;
		1771: SAMPLE = 16'h34c4;
		1772: SAMPLE = 16'h3496;
		1773: SAMPLE = 16'h3468;
		1774: SAMPLE = 16'h343a;
		1775: SAMPLE = 16'h340c;
		1776: SAMPLE = 16'h33de;
		1777: SAMPLE = 16'h33b0;
		1778: SAMPLE = 16'h3382;
		1779: SAMPLE = 16'h3354;
		1780: SAMPLE = 16'h3326;
		1781: SAMPLE = 16'h32f8;
		1782: SAMPLE = 16'h32ca;
		1783: SAMPLE = 16'h329c;
		1784: SAMPLE = 16'h326e;
		1785: SAMPLE = 16'h3240;
		1786: SAMPLE = 16'h3211;
		1787: SAMPLE = 16'h31e3;
		1788: SAMPLE = 16'h31b5;
		1789: SAMPLE = 16'h3186;
		1790: SAMPLE = 16'h3158;
		1791: SAMPLE = 16'h312a;
		1792: SAMPLE = 16'h30fb;
		1793: SAMPLE = 16'h30cd;
		1794: SAMPLE = 16'h309e;
		1795: SAMPLE = 16'h3070;
		1796: SAMPLE = 16'h3041;
		1797: SAMPLE = 16'h3013;
		1798: SAMPLE = 16'h2fe4;
		1799: SAMPLE = 16'h2fb5;
		1800: SAMPLE = 16'h2f87;
		1801: SAMPLE = 16'h2f58;
		1802: SAMPLE = 16'h2f29;
		1803: SAMPLE = 16'h2efb;
		1804: SAMPLE = 16'h2ecc;
		1805: SAMPLE = 16'h2e9d;
		1806: SAMPLE = 16'h2e6e;
		1807: SAMPLE = 16'h2e3f;
		1808: SAMPLE = 16'h2e11;
		1809: SAMPLE = 16'h2de2;
		1810: SAMPLE = 16'h2db3;
		1811: SAMPLE = 16'h2d84;
		1812: SAMPLE = 16'h2d55;
		1813: SAMPLE = 16'h2d26;
		1814: SAMPLE = 16'h2cf7;
		1815: SAMPLE = 16'h2cc8;
		1816: SAMPLE = 16'h2c98;
		1817: SAMPLE = 16'h2c69;
		1818: SAMPLE = 16'h2c3a;
		1819: SAMPLE = 16'h2c0b;
		1820: SAMPLE = 16'h2bdc;
		1821: SAMPLE = 16'h2bad;
		1822: SAMPLE = 16'h2b7d;
		1823: SAMPLE = 16'h2b4e;
		1824: SAMPLE = 16'h2b1f;
		1825: SAMPLE = 16'h2aef;
		1826: SAMPLE = 16'h2ac0;
		1827: SAMPLE = 16'h2a91;
		1828: SAMPLE = 16'h2a61;
		1829: SAMPLE = 16'h2a32;
		1830: SAMPLE = 16'h2a02;
		1831: SAMPLE = 16'h29d3;
		1832: SAMPLE = 16'h29a3;
		1833: SAMPLE = 16'h2974;
		1834: SAMPLE = 16'h2944;
		1835: SAMPLE = 16'h2915;
		1836: SAMPLE = 16'h28e5;
		1837: SAMPLE = 16'h28b5;
		1838: SAMPLE = 16'h2886;
		1839: SAMPLE = 16'h2856;
		1840: SAMPLE = 16'h2826;
		1841: SAMPLE = 16'h27f6;
		1842: SAMPLE = 16'h27c7;
		1843: SAMPLE = 16'h2797;
		1844: SAMPLE = 16'h2767;
		1845: SAMPLE = 16'h2737;
		1846: SAMPLE = 16'h2707;
		1847: SAMPLE = 16'h26d8;
		1848: SAMPLE = 16'h26a8;
		1849: SAMPLE = 16'h2678;
		1850: SAMPLE = 16'h2648;
		1851: SAMPLE = 16'h2618;
		1852: SAMPLE = 16'h25e8;
		1853: SAMPLE = 16'h25b8;
		1854: SAMPLE = 16'h2588;
		1855: SAMPLE = 16'h2558;
		1856: SAMPLE = 16'h2528;
		1857: SAMPLE = 16'h24f7;
		1858: SAMPLE = 16'h24c7;
		1859: SAMPLE = 16'h2497;
		1860: SAMPLE = 16'h2467;
		1861: SAMPLE = 16'h2437;
		1862: SAMPLE = 16'h2407;
		1863: SAMPLE = 16'h23d6;
		1864: SAMPLE = 16'h23a6;
		1865: SAMPLE = 16'h2376;
		1866: SAMPLE = 16'h2345;
		1867: SAMPLE = 16'h2315;
		1868: SAMPLE = 16'h22e5;
		1869: SAMPLE = 16'h22b4;
		1870: SAMPLE = 16'h2284;
		1871: SAMPLE = 16'h2254;
		1872: SAMPLE = 16'h2223;
		1873: SAMPLE = 16'h21f3;
		1874: SAMPLE = 16'h21c2;
		1875: SAMPLE = 16'h2192;
		1876: SAMPLE = 16'h2161;
		1877: SAMPLE = 16'h2131;
		1878: SAMPLE = 16'h2100;
		1879: SAMPLE = 16'h20d0;
		1880: SAMPLE = 16'h209f;
		1881: SAMPLE = 16'h206e;
		1882: SAMPLE = 16'h203e;
		1883: SAMPLE = 16'h200d;
		1884: SAMPLE = 16'h1fdc;
		1885: SAMPLE = 16'h1fac;
		1886: SAMPLE = 16'h1f7b;
		1887: SAMPLE = 16'h1f4a;
		1888: SAMPLE = 16'h1f19;
		1889: SAMPLE = 16'h1ee9;
		1890: SAMPLE = 16'h1eb8;
		1891: SAMPLE = 16'h1e87;
		1892: SAMPLE = 16'h1e56;
		1893: SAMPLE = 16'h1e25;
		1894: SAMPLE = 16'h1df5;
		1895: SAMPLE = 16'h1dc4;
		1896: SAMPLE = 16'h1d93;
		1897: SAMPLE = 16'h1d62;
		1898: SAMPLE = 16'h1d31;
		1899: SAMPLE = 16'h1d00;
		1900: SAMPLE = 16'h1ccf;
		1901: SAMPLE = 16'h1c9e;
		1902: SAMPLE = 16'h1c6d;
		1903: SAMPLE = 16'h1c3c;
		1904: SAMPLE = 16'h1c0b;
		1905: SAMPLE = 16'h1bda;
		1906: SAMPLE = 16'h1ba9;
		1907: SAMPLE = 16'h1b78;
		1908: SAMPLE = 16'h1b47;
		1909: SAMPLE = 16'h1b16;
		1910: SAMPLE = 16'h1ae4;
		1911: SAMPLE = 16'h1ab3;
		1912: SAMPLE = 16'h1a82;
		1913: SAMPLE = 16'h1a51;
		1914: SAMPLE = 16'h1a20;
		1915: SAMPLE = 16'h19ef;
		1916: SAMPLE = 16'h19bd;
		1917: SAMPLE = 16'h198c;
		1918: SAMPLE = 16'h195b;
		1919: SAMPLE = 16'h192a;
		1920: SAMPLE = 16'h18f8;
		1921: SAMPLE = 16'h18c7;
		1922: SAMPLE = 16'h1896;
		1923: SAMPLE = 16'h1864;
		1924: SAMPLE = 16'h1833;
		1925: SAMPLE = 16'h1802;
		1926: SAMPLE = 16'h17d0;
		1927: SAMPLE = 16'h179f;
		1928: SAMPLE = 16'h176d;
		1929: SAMPLE = 16'h173c;
		1930: SAMPLE = 16'h170a;
		1931: SAMPLE = 16'h16d9;
		1932: SAMPLE = 16'h16a8;
		1933: SAMPLE = 16'h1676;
		1934: SAMPLE = 16'h1645;
		1935: SAMPLE = 16'h1613;
		1936: SAMPLE = 16'h15e2;
		1937: SAMPLE = 16'h15b0;
		1938: SAMPLE = 16'h157f;
		1939: SAMPLE = 16'h154d;
		1940: SAMPLE = 16'h151b;
		1941: SAMPLE = 16'h14ea;
		1942: SAMPLE = 16'h14b8;
		1943: SAMPLE = 16'h1487;
		1944: SAMPLE = 16'h1455;
		1945: SAMPLE = 16'h1423;
		1946: SAMPLE = 16'h13f2;
		1947: SAMPLE = 16'h13c0;
		1948: SAMPLE = 16'h138e;
		1949: SAMPLE = 16'h135d;
		1950: SAMPLE = 16'h132b;
		1951: SAMPLE = 16'h12f9;
		1952: SAMPLE = 16'h12c8;
		1953: SAMPLE = 16'h1296;
		1954: SAMPLE = 16'h1264;
		1955: SAMPLE = 16'h1232;
		1956: SAMPLE = 16'h1201;
		1957: SAMPLE = 16'h11cf;
		1958: SAMPLE = 16'h119d;
		1959: SAMPLE = 16'h116b;
		1960: SAMPLE = 16'h1139;
		1961: SAMPLE = 16'h1108;
		1962: SAMPLE = 16'h10d6;
		1963: SAMPLE = 16'h10a4;
		1964: SAMPLE = 16'h1072;
		1965: SAMPLE = 16'h1040;
		1966: SAMPLE = 16'h100e;
		1967: SAMPLE = 16'hfdd;
		1968: SAMPLE = 16'hfab;
		1969: SAMPLE = 16'hf79;
		1970: SAMPLE = 16'hf47;
		1971: SAMPLE = 16'hf15;
		1972: SAMPLE = 16'hee3;
		1973: SAMPLE = 16'heb1;
		1974: SAMPLE = 16'he7f;
		1975: SAMPLE = 16'he4d;
		1976: SAMPLE = 16'he1b;
		1977: SAMPLE = 16'hde9;
		1978: SAMPLE = 16'hdb7;
		1979: SAMPLE = 16'hd85;
		1980: SAMPLE = 16'hd53;
		1981: SAMPLE = 16'hd21;
		1982: SAMPLE = 16'hcef;
		1983: SAMPLE = 16'hcbd;
		1984: SAMPLE = 16'hc8b;
		1985: SAMPLE = 16'hc59;
		1986: SAMPLE = 16'hc27;
		1987: SAMPLE = 16'hbf5;
		1988: SAMPLE = 16'hbc3;
		1989: SAMPLE = 16'hb91;
		1990: SAMPLE = 16'hb5f;
		1991: SAMPLE = 16'hb2d;
		1992: SAMPLE = 16'hafb;
		1993: SAMPLE = 16'hac9;
		1994: SAMPLE = 16'ha97;
		1995: SAMPLE = 16'ha65;
		1996: SAMPLE = 16'ha33;
		1997: SAMPLE = 16'ha00;
		1998: SAMPLE = 16'h9ce;
		1999: SAMPLE = 16'h99c;
		2000: SAMPLE = 16'h96a;
		2001: SAMPLE = 16'h938;
		2002: SAMPLE = 16'h906;
		2003: SAMPLE = 16'h8d4;
		2004: SAMPLE = 16'h8a2;
		2005: SAMPLE = 16'h86f;
		2006: SAMPLE = 16'h83d;
		2007: SAMPLE = 16'h80b;
		2008: SAMPLE = 16'h7d9;
		2009: SAMPLE = 16'h7a7;
		2010: SAMPLE = 16'h775;
		2011: SAMPLE = 16'h742;
		2012: SAMPLE = 16'h710;
		2013: SAMPLE = 16'h6de;
		2014: SAMPLE = 16'h6ac;
		2015: SAMPLE = 16'h67a;
		2016: SAMPLE = 16'h647;
		2017: SAMPLE = 16'h615;
		2018: SAMPLE = 16'h5e3;
		2019: SAMPLE = 16'h5b1;
		2020: SAMPLE = 16'h57f;
		2021: SAMPLE = 16'h54c;
		2022: SAMPLE = 16'h51a;
		2023: SAMPLE = 16'h4e8;
		2024: SAMPLE = 16'h4b6;
		2025: SAMPLE = 16'h483;
		2026: SAMPLE = 16'h451;
		2027: SAMPLE = 16'h41f;
		2028: SAMPLE = 16'h3ed;
		2029: SAMPLE = 16'h3ba;
		2030: SAMPLE = 16'h388;
		2031: SAMPLE = 16'h356;
		2032: SAMPLE = 16'h324;
		2033: SAMPLE = 16'h2f1;
		2034: SAMPLE = 16'h2bf;
		2035: SAMPLE = 16'h28d;
		2036: SAMPLE = 16'h25b;
		2037: SAMPLE = 16'h228;
		2038: SAMPLE = 16'h1f6;
		2039: SAMPLE = 16'h1c4;
		2040: SAMPLE = 16'h192;
		2041: SAMPLE = 16'h15f;
		2042: SAMPLE = 16'h12d;
		2043: SAMPLE = 16'hfb;
		2044: SAMPLE = 16'hc9;
		2045: SAMPLE = 16'h96;
		2046: SAMPLE = 16'h64;
		2047: SAMPLE = 16'h32;
		2048: SAMPLE = 16'h0;
		2049: SAMPLE = 16'hffcd;
		2050: SAMPLE = 16'hff9b;
		2051: SAMPLE = 16'hff69;
		2052: SAMPLE = 16'hff36;
		2053: SAMPLE = 16'hff04;
		2054: SAMPLE = 16'hfed2;
		2055: SAMPLE = 16'hfea0;
		2056: SAMPLE = 16'hfe6d;
		2057: SAMPLE = 16'hfe3b;
		2058: SAMPLE = 16'hfe09;
		2059: SAMPLE = 16'hfdd7;
		2060: SAMPLE = 16'hfda4;
		2061: SAMPLE = 16'hfd72;
		2062: SAMPLE = 16'hfd40;
		2063: SAMPLE = 16'hfd0e;
		2064: SAMPLE = 16'hfcdb;
		2065: SAMPLE = 16'hfca9;
		2066: SAMPLE = 16'hfc77;
		2067: SAMPLE = 16'hfc45;
		2068: SAMPLE = 16'hfc12;
		2069: SAMPLE = 16'hfbe0;
		2070: SAMPLE = 16'hfbae;
		2071: SAMPLE = 16'hfb7c;
		2072: SAMPLE = 16'hfb49;
		2073: SAMPLE = 16'hfb17;
		2074: SAMPLE = 16'hfae5;
		2075: SAMPLE = 16'hfab3;
		2076: SAMPLE = 16'hfa80;
		2077: SAMPLE = 16'hfa4e;
		2078: SAMPLE = 16'hfa1c;
		2079: SAMPLE = 16'hf9ea;
		2080: SAMPLE = 16'hf9b8;
		2081: SAMPLE = 16'hf985;
		2082: SAMPLE = 16'hf953;
		2083: SAMPLE = 16'hf921;
		2084: SAMPLE = 16'hf8ef;
		2085: SAMPLE = 16'hf8bd;
		2086: SAMPLE = 16'hf88a;
		2087: SAMPLE = 16'hf858;
		2088: SAMPLE = 16'hf826;
		2089: SAMPLE = 16'hf7f4;
		2090: SAMPLE = 16'hf7c2;
		2091: SAMPLE = 16'hf790;
		2092: SAMPLE = 16'hf75d;
		2093: SAMPLE = 16'hf72b;
		2094: SAMPLE = 16'hf6f9;
		2095: SAMPLE = 16'hf6c7;
		2096: SAMPLE = 16'hf695;
		2097: SAMPLE = 16'hf663;
		2098: SAMPLE = 16'hf631;
		2099: SAMPLE = 16'hf5ff;
		2100: SAMPLE = 16'hf5cc;
		2101: SAMPLE = 16'hf59a;
		2102: SAMPLE = 16'hf568;
		2103: SAMPLE = 16'hf536;
		2104: SAMPLE = 16'hf504;
		2105: SAMPLE = 16'hf4d2;
		2106: SAMPLE = 16'hf4a0;
		2107: SAMPLE = 16'hf46e;
		2108: SAMPLE = 16'hf43c;
		2109: SAMPLE = 16'hf40a;
		2110: SAMPLE = 16'hf3d8;
		2111: SAMPLE = 16'hf3a6;
		2112: SAMPLE = 16'hf374;
		2113: SAMPLE = 16'hf342;
		2114: SAMPLE = 16'hf310;
		2115: SAMPLE = 16'hf2de;
		2116: SAMPLE = 16'hf2ac;
		2117: SAMPLE = 16'hf27a;
		2118: SAMPLE = 16'hf248;
		2119: SAMPLE = 16'hf216;
		2120: SAMPLE = 16'hf1e4;
		2121: SAMPLE = 16'hf1b2;
		2122: SAMPLE = 16'hf180;
		2123: SAMPLE = 16'hf14e;
		2124: SAMPLE = 16'hf11c;
		2125: SAMPLE = 16'hf0ea;
		2126: SAMPLE = 16'hf0b8;
		2127: SAMPLE = 16'hf086;
		2128: SAMPLE = 16'hf054;
		2129: SAMPLE = 16'hf022;
		2130: SAMPLE = 16'heff1;
		2131: SAMPLE = 16'hefbf;
		2132: SAMPLE = 16'hef8d;
		2133: SAMPLE = 16'hef5b;
		2134: SAMPLE = 16'hef29;
		2135: SAMPLE = 16'heef7;
		2136: SAMPLE = 16'heec6;
		2137: SAMPLE = 16'hee94;
		2138: SAMPLE = 16'hee62;
		2139: SAMPLE = 16'hee30;
		2140: SAMPLE = 16'hedfe;
		2141: SAMPLE = 16'hedcd;
		2142: SAMPLE = 16'hed9b;
		2143: SAMPLE = 16'hed69;
		2144: SAMPLE = 16'hed37;
		2145: SAMPLE = 16'hed06;
		2146: SAMPLE = 16'hecd4;
		2147: SAMPLE = 16'heca2;
		2148: SAMPLE = 16'hec71;
		2149: SAMPLE = 16'hec3f;
		2150: SAMPLE = 16'hec0d;
		2151: SAMPLE = 16'hebdc;
		2152: SAMPLE = 16'hebaa;
		2153: SAMPLE = 16'heb78;
		2154: SAMPLE = 16'heb47;
		2155: SAMPLE = 16'heb15;
		2156: SAMPLE = 16'heae4;
		2157: SAMPLE = 16'heab2;
		2158: SAMPLE = 16'hea80;
		2159: SAMPLE = 16'hea4f;
		2160: SAMPLE = 16'hea1d;
		2161: SAMPLE = 16'he9ec;
		2162: SAMPLE = 16'he9ba;
		2163: SAMPLE = 16'he989;
		2164: SAMPLE = 16'he957;
		2165: SAMPLE = 16'he926;
		2166: SAMPLE = 16'he8f5;
		2167: SAMPLE = 16'he8c3;
		2168: SAMPLE = 16'he892;
		2169: SAMPLE = 16'he860;
		2170: SAMPLE = 16'he82f;
		2171: SAMPLE = 16'he7fd;
		2172: SAMPLE = 16'he7cc;
		2173: SAMPLE = 16'he79b;
		2174: SAMPLE = 16'he769;
		2175: SAMPLE = 16'he738;
		2176: SAMPLE = 16'he707;
		2177: SAMPLE = 16'he6d5;
		2178: SAMPLE = 16'he6a4;
		2179: SAMPLE = 16'he673;
		2180: SAMPLE = 16'he642;
		2181: SAMPLE = 16'he610;
		2182: SAMPLE = 16'he5df;
		2183: SAMPLE = 16'he5ae;
		2184: SAMPLE = 16'he57d;
		2185: SAMPLE = 16'he54c;
		2186: SAMPLE = 16'he51b;
		2187: SAMPLE = 16'he4e9;
		2188: SAMPLE = 16'he4b8;
		2189: SAMPLE = 16'he487;
		2190: SAMPLE = 16'he456;
		2191: SAMPLE = 16'he425;
		2192: SAMPLE = 16'he3f4;
		2193: SAMPLE = 16'he3c3;
		2194: SAMPLE = 16'he392;
		2195: SAMPLE = 16'he361;
		2196: SAMPLE = 16'he330;
		2197: SAMPLE = 16'he2ff;
		2198: SAMPLE = 16'he2ce;
		2199: SAMPLE = 16'he29d;
		2200: SAMPLE = 16'he26c;
		2201: SAMPLE = 16'he23b;
		2202: SAMPLE = 16'he20a;
		2203: SAMPLE = 16'he1da;
		2204: SAMPLE = 16'he1a9;
		2205: SAMPLE = 16'he178;
		2206: SAMPLE = 16'he147;
		2207: SAMPLE = 16'he116;
		2208: SAMPLE = 16'he0e6;
		2209: SAMPLE = 16'he0b5;
		2210: SAMPLE = 16'he084;
		2211: SAMPLE = 16'he053;
		2212: SAMPLE = 16'he023;
		2213: SAMPLE = 16'hdff2;
		2214: SAMPLE = 16'hdfc1;
		2215: SAMPLE = 16'hdf91;
		2216: SAMPLE = 16'hdf60;
		2217: SAMPLE = 16'hdf2f;
		2218: SAMPLE = 16'hdeff;
		2219: SAMPLE = 16'hdece;
		2220: SAMPLE = 16'hde9e;
		2221: SAMPLE = 16'hde6d;
		2222: SAMPLE = 16'hde3d;
		2223: SAMPLE = 16'hde0c;
		2224: SAMPLE = 16'hdddc;
		2225: SAMPLE = 16'hddab;
		2226: SAMPLE = 16'hdd7b;
		2227: SAMPLE = 16'hdd4b;
		2228: SAMPLE = 16'hdd1a;
		2229: SAMPLE = 16'hdcea;
		2230: SAMPLE = 16'hdcba;
		2231: SAMPLE = 16'hdc89;
		2232: SAMPLE = 16'hdc59;
		2233: SAMPLE = 16'hdc29;
		2234: SAMPLE = 16'hdbf8;
		2235: SAMPLE = 16'hdbc8;
		2236: SAMPLE = 16'hdb98;
		2237: SAMPLE = 16'hdb68;
		2238: SAMPLE = 16'hdb38;
		2239: SAMPLE = 16'hdb08;
		2240: SAMPLE = 16'hdad7;
		2241: SAMPLE = 16'hdaa7;
		2242: SAMPLE = 16'hda77;
		2243: SAMPLE = 16'hda47;
		2244: SAMPLE = 16'hda17;
		2245: SAMPLE = 16'hd9e7;
		2246: SAMPLE = 16'hd9b7;
		2247: SAMPLE = 16'hd987;
		2248: SAMPLE = 16'hd957;
		2249: SAMPLE = 16'hd927;
		2250: SAMPLE = 16'hd8f8;
		2251: SAMPLE = 16'hd8c8;
		2252: SAMPLE = 16'hd898;
		2253: SAMPLE = 16'hd868;
		2254: SAMPLE = 16'hd838;
		2255: SAMPLE = 16'hd809;
		2256: SAMPLE = 16'hd7d9;
		2257: SAMPLE = 16'hd7a9;
		2258: SAMPLE = 16'hd779;
		2259: SAMPLE = 16'hd74a;
		2260: SAMPLE = 16'hd71a;
		2261: SAMPLE = 16'hd6ea;
		2262: SAMPLE = 16'hd6bb;
		2263: SAMPLE = 16'hd68b;
		2264: SAMPLE = 16'hd65c;
		2265: SAMPLE = 16'hd62c;
		2266: SAMPLE = 16'hd5fd;
		2267: SAMPLE = 16'hd5cd;
		2268: SAMPLE = 16'hd59e;
		2269: SAMPLE = 16'hd56e;
		2270: SAMPLE = 16'hd53f;
		2271: SAMPLE = 16'hd510;
		2272: SAMPLE = 16'hd4e0;
		2273: SAMPLE = 16'hd4b1;
		2274: SAMPLE = 16'hd482;
		2275: SAMPLE = 16'hd452;
		2276: SAMPLE = 16'hd423;
		2277: SAMPLE = 16'hd3f4;
		2278: SAMPLE = 16'hd3c5;
		2279: SAMPLE = 16'hd396;
		2280: SAMPLE = 16'hd367;
		2281: SAMPLE = 16'hd337;
		2282: SAMPLE = 16'hd308;
		2283: SAMPLE = 16'hd2d9;
		2284: SAMPLE = 16'hd2aa;
		2285: SAMPLE = 16'hd27b;
		2286: SAMPLE = 16'hd24c;
		2287: SAMPLE = 16'hd21d;
		2288: SAMPLE = 16'hd1ee;
		2289: SAMPLE = 16'hd1c0;
		2290: SAMPLE = 16'hd191;
		2291: SAMPLE = 16'hd162;
		2292: SAMPLE = 16'hd133;
		2293: SAMPLE = 16'hd104;
		2294: SAMPLE = 16'hd0d6;
		2295: SAMPLE = 16'hd0a7;
		2296: SAMPLE = 16'hd078;
		2297: SAMPLE = 16'hd04a;
		2298: SAMPLE = 16'hd01b;
		2299: SAMPLE = 16'hcfec;
		2300: SAMPLE = 16'hcfbe;
		2301: SAMPLE = 16'hcf8f;
		2302: SAMPLE = 16'hcf61;
		2303: SAMPLE = 16'hcf32;
		2304: SAMPLE = 16'hcf04;
		2305: SAMPLE = 16'hced5;
		2306: SAMPLE = 16'hcea7;
		2307: SAMPLE = 16'hce79;
		2308: SAMPLE = 16'hce4a;
		2309: SAMPLE = 16'hce1c;
		2310: SAMPLE = 16'hcdee;
		2311: SAMPLE = 16'hcdbf;
		2312: SAMPLE = 16'hcd91;
		2313: SAMPLE = 16'hcd63;
		2314: SAMPLE = 16'hcd35;
		2315: SAMPLE = 16'hcd07;
		2316: SAMPLE = 16'hccd9;
		2317: SAMPLE = 16'hccab;
		2318: SAMPLE = 16'hcc7d;
		2319: SAMPLE = 16'hcc4f;
		2320: SAMPLE = 16'hcc21;
		2321: SAMPLE = 16'hcbf3;
		2322: SAMPLE = 16'hcbc5;
		2323: SAMPLE = 16'hcb97;
		2324: SAMPLE = 16'hcb69;
		2325: SAMPLE = 16'hcb3b;
		2326: SAMPLE = 16'hcb0d;
		2327: SAMPLE = 16'hcae0;
		2328: SAMPLE = 16'hcab2;
		2329: SAMPLE = 16'hca84;
		2330: SAMPLE = 16'hca57;
		2331: SAMPLE = 16'hca29;
		2332: SAMPLE = 16'hc9fb;
		2333: SAMPLE = 16'hc9ce;
		2334: SAMPLE = 16'hc9a0;
		2335: SAMPLE = 16'hc973;
		2336: SAMPLE = 16'hc945;
		2337: SAMPLE = 16'hc918;
		2338: SAMPLE = 16'hc8eb;
		2339: SAMPLE = 16'hc8bd;
		2340: SAMPLE = 16'hc890;
		2341: SAMPLE = 16'hc863;
		2342: SAMPLE = 16'hc835;
		2343: SAMPLE = 16'hc808;
		2344: SAMPLE = 16'hc7db;
		2345: SAMPLE = 16'hc7ae;
		2346: SAMPLE = 16'hc781;
		2347: SAMPLE = 16'hc754;
		2348: SAMPLE = 16'hc727;
		2349: SAMPLE = 16'hc6f9;
		2350: SAMPLE = 16'hc6cd;
		2351: SAMPLE = 16'hc6a0;
		2352: SAMPLE = 16'hc673;
		2353: SAMPLE = 16'hc646;
		2354: SAMPLE = 16'hc619;
		2355: SAMPLE = 16'hc5ec;
		2356: SAMPLE = 16'hc5bf;
		2357: SAMPLE = 16'hc593;
		2358: SAMPLE = 16'hc566;
		2359: SAMPLE = 16'hc539;
		2360: SAMPLE = 16'hc50d;
		2361: SAMPLE = 16'hc4e0;
		2362: SAMPLE = 16'hc4b3;
		2363: SAMPLE = 16'hc487;
		2364: SAMPLE = 16'hc45a;
		2365: SAMPLE = 16'hc42e;
		2366: SAMPLE = 16'hc402;
		2367: SAMPLE = 16'hc3d5;
		2368: SAMPLE = 16'hc3a9;
		2369: SAMPLE = 16'hc37c;
		2370: SAMPLE = 16'hc350;
		2371: SAMPLE = 16'hc324;
		2372: SAMPLE = 16'hc2f8;
		2373: SAMPLE = 16'hc2cc;
		2374: SAMPLE = 16'hc29f;
		2375: SAMPLE = 16'hc273;
		2376: SAMPLE = 16'hc247;
		2377: SAMPLE = 16'hc21b;
		2378: SAMPLE = 16'hc1ef;
		2379: SAMPLE = 16'hc1c3;
		2380: SAMPLE = 16'hc197;
		2381: SAMPLE = 16'hc16c;
		2382: SAMPLE = 16'hc140;
		2383: SAMPLE = 16'hc114;
		2384: SAMPLE = 16'hc0e8;
		2385: SAMPLE = 16'hc0bc;
		2386: SAMPLE = 16'hc091;
		2387: SAMPLE = 16'hc065;
		2388: SAMPLE = 16'hc03a;
		2389: SAMPLE = 16'hc00e;
		2390: SAMPLE = 16'hbfe2;
		2391: SAMPLE = 16'hbfb7;
		2392: SAMPLE = 16'hbf8c;
		2393: SAMPLE = 16'hbf60;
		2394: SAMPLE = 16'hbf35;
		2395: SAMPLE = 16'hbf09;
		2396: SAMPLE = 16'hbede;
		2397: SAMPLE = 16'hbeb3;
		2398: SAMPLE = 16'hbe88;
		2399: SAMPLE = 16'hbe5d;
		2400: SAMPLE = 16'hbe31;
		2401: SAMPLE = 16'hbe06;
		2402: SAMPLE = 16'hbddb;
		2403: SAMPLE = 16'hbdb0;
		2404: SAMPLE = 16'hbd85;
		2405: SAMPLE = 16'hbd5a;
		2406: SAMPLE = 16'hbd2f;
		2407: SAMPLE = 16'hbd05;
		2408: SAMPLE = 16'hbcda;
		2409: SAMPLE = 16'hbcaf;
		2410: SAMPLE = 16'hbc84;
		2411: SAMPLE = 16'hbc5a;
		2412: SAMPLE = 16'hbc2f;
		2413: SAMPLE = 16'hbc04;
		2414: SAMPLE = 16'hbbda;
		2415: SAMPLE = 16'hbbaf;
		2416: SAMPLE = 16'hbb85;
		2417: SAMPLE = 16'hbb5a;
		2418: SAMPLE = 16'hbb30;
		2419: SAMPLE = 16'hbb05;
		2420: SAMPLE = 16'hbadb;
		2421: SAMPLE = 16'hbab1;
		2422: SAMPLE = 16'hba87;
		2423: SAMPLE = 16'hba5c;
		2424: SAMPLE = 16'hba32;
		2425: SAMPLE = 16'hba08;
		2426: SAMPLE = 16'hb9de;
		2427: SAMPLE = 16'hb9b4;
		2428: SAMPLE = 16'hb98a;
		2429: SAMPLE = 16'hb960;
		2430: SAMPLE = 16'hb936;
		2431: SAMPLE = 16'hb90c;
		2432: SAMPLE = 16'hb8e3;
		2433: SAMPLE = 16'hb8b9;
		2434: SAMPLE = 16'hb88f;
		2435: SAMPLE = 16'hb865;
		2436: SAMPLE = 16'hb83c;
		2437: SAMPLE = 16'hb812;
		2438: SAMPLE = 16'hb7e9;
		2439: SAMPLE = 16'hb7bf;
		2440: SAMPLE = 16'hb796;
		2441: SAMPLE = 16'hb76c;
		2442: SAMPLE = 16'hb743;
		2443: SAMPLE = 16'hb719;
		2444: SAMPLE = 16'hb6f0;
		2445: SAMPLE = 16'hb6c7;
		2446: SAMPLE = 16'hb69e;
		2447: SAMPLE = 16'hb675;
		2448: SAMPLE = 16'hb64b;
		2449: SAMPLE = 16'hb622;
		2450: SAMPLE = 16'hb5f9;
		2451: SAMPLE = 16'hb5d0;
		2452: SAMPLE = 16'hb5a7;
		2453: SAMPLE = 16'hb57e;
		2454: SAMPLE = 16'hb556;
		2455: SAMPLE = 16'hb52d;
		2456: SAMPLE = 16'hb504;
		2457: SAMPLE = 16'hb4db;
		2458: SAMPLE = 16'hb4b3;
		2459: SAMPLE = 16'hb48a;
		2460: SAMPLE = 16'hb461;
		2461: SAMPLE = 16'hb439;
		2462: SAMPLE = 16'hb410;
		2463: SAMPLE = 16'hb3e8;
		2464: SAMPLE = 16'hb3c0;
		2465: SAMPLE = 16'hb397;
		2466: SAMPLE = 16'hb36f;
		2467: SAMPLE = 16'hb347;
		2468: SAMPLE = 16'hb31e;
		2469: SAMPLE = 16'hb2f6;
		2470: SAMPLE = 16'hb2ce;
		2471: SAMPLE = 16'hb2a6;
		2472: SAMPLE = 16'hb27e;
		2473: SAMPLE = 16'hb256;
		2474: SAMPLE = 16'hb22e;
		2475: SAMPLE = 16'hb206;
		2476: SAMPLE = 16'hb1de;
		2477: SAMPLE = 16'hb1b7;
		2478: SAMPLE = 16'hb18f;
		2479: SAMPLE = 16'hb167;
		2480: SAMPLE = 16'hb140;
		2481: SAMPLE = 16'hb118;
		2482: SAMPLE = 16'hb0f0;
		2483: SAMPLE = 16'hb0c9;
		2484: SAMPLE = 16'hb0a1;
		2485: SAMPLE = 16'hb07a;
		2486: SAMPLE = 16'hb053;
		2487: SAMPLE = 16'hb02b;
		2488: SAMPLE = 16'hb004;
		2489: SAMPLE = 16'hafdd;
		2490: SAMPLE = 16'hafb6;
		2491: SAMPLE = 16'haf8f;
		2492: SAMPLE = 16'haf68;
		2493: SAMPLE = 16'haf40;
		2494: SAMPLE = 16'haf1a;
		2495: SAMPLE = 16'haef3;
		2496: SAMPLE = 16'haecc;
		2497: SAMPLE = 16'haea5;
		2498: SAMPLE = 16'hae7e;
		2499: SAMPLE = 16'hae57;
		2500: SAMPLE = 16'hae31;
		2501: SAMPLE = 16'hae0a;
		2502: SAMPLE = 16'hade3;
		2503: SAMPLE = 16'hadbd;
		2504: SAMPLE = 16'had96;
		2505: SAMPLE = 16'had70;
		2506: SAMPLE = 16'had4a;
		2507: SAMPLE = 16'had23;
		2508: SAMPLE = 16'hacfd;
		2509: SAMPLE = 16'hacd7;
		2510: SAMPLE = 16'hacb1;
		2511: SAMPLE = 16'hac8a;
		2512: SAMPLE = 16'hac64;
		2513: SAMPLE = 16'hac3e;
		2514: SAMPLE = 16'hac18;
		2515: SAMPLE = 16'habf2;
		2516: SAMPLE = 16'habcc;
		2517: SAMPLE = 16'haba7;
		2518: SAMPLE = 16'hab81;
		2519: SAMPLE = 16'hab5b;
		2520: SAMPLE = 16'hab35;
		2521: SAMPLE = 16'hab10;
		2522: SAMPLE = 16'haaea;
		2523: SAMPLE = 16'haac5;
		2524: SAMPLE = 16'haa9f;
		2525: SAMPLE = 16'haa7a;
		2526: SAMPLE = 16'haa54;
		2527: SAMPLE = 16'haa2f;
		2528: SAMPLE = 16'haa0a;
		2529: SAMPLE = 16'ha9e5;
		2530: SAMPLE = 16'ha9bf;
		2531: SAMPLE = 16'ha99a;
		2532: SAMPLE = 16'ha975;
		2533: SAMPLE = 16'ha950;
		2534: SAMPLE = 16'ha92b;
		2535: SAMPLE = 16'ha906;
		2536: SAMPLE = 16'ha8e2;
		2537: SAMPLE = 16'ha8bd;
		2538: SAMPLE = 16'ha898;
		2539: SAMPLE = 16'ha873;
		2540: SAMPLE = 16'ha84f;
		2541: SAMPLE = 16'ha82a;
		2542: SAMPLE = 16'ha806;
		2543: SAMPLE = 16'ha7e1;
		2544: SAMPLE = 16'ha7bd;
		2545: SAMPLE = 16'ha798;
		2546: SAMPLE = 16'ha774;
		2547: SAMPLE = 16'ha750;
		2548: SAMPLE = 16'ha72b;
		2549: SAMPLE = 16'ha707;
		2550: SAMPLE = 16'ha6e3;
		2551: SAMPLE = 16'ha6bf;
		2552: SAMPLE = 16'ha69b;
		2553: SAMPLE = 16'ha677;
		2554: SAMPLE = 16'ha653;
		2555: SAMPLE = 16'ha62f;
		2556: SAMPLE = 16'ha60c;
		2557: SAMPLE = 16'ha5e8;
		2558: SAMPLE = 16'ha5c4;
		2559: SAMPLE = 16'ha5a1;
		2560: SAMPLE = 16'ha57d;
		2561: SAMPLE = 16'ha55a;
		2562: SAMPLE = 16'ha536;
		2563: SAMPLE = 16'ha513;
		2564: SAMPLE = 16'ha4ef;
		2565: SAMPLE = 16'ha4cc;
		2566: SAMPLE = 16'ha4a9;
		2567: SAMPLE = 16'ha486;
		2568: SAMPLE = 16'ha462;
		2569: SAMPLE = 16'ha43f;
		2570: SAMPLE = 16'ha41c;
		2571: SAMPLE = 16'ha3f9;
		2572: SAMPLE = 16'ha3d6;
		2573: SAMPLE = 16'ha3b4;
		2574: SAMPLE = 16'ha391;
		2575: SAMPLE = 16'ha36e;
		2576: SAMPLE = 16'ha34b;
		2577: SAMPLE = 16'ha329;
		2578: SAMPLE = 16'ha306;
		2579: SAMPLE = 16'ha2e4;
		2580: SAMPLE = 16'ha2c1;
		2581: SAMPLE = 16'ha29f;
		2582: SAMPLE = 16'ha27c;
		2583: SAMPLE = 16'ha25a;
		2584: SAMPLE = 16'ha238;
		2585: SAMPLE = 16'ha216;
		2586: SAMPLE = 16'ha1f4;
		2587: SAMPLE = 16'ha1d2;
		2588: SAMPLE = 16'ha1af;
		2589: SAMPLE = 16'ha18e;
		2590: SAMPLE = 16'ha16c;
		2591: SAMPLE = 16'ha14a;
		2592: SAMPLE = 16'ha128;
		2593: SAMPLE = 16'ha106;
		2594: SAMPLE = 16'ha0e5;
		2595: SAMPLE = 16'ha0c3;
		2596: SAMPLE = 16'ha0a1;
		2597: SAMPLE = 16'ha080;
		2598: SAMPLE = 16'ha05f;
		2599: SAMPLE = 16'ha03d;
		2600: SAMPLE = 16'ha01c;
		2601: SAMPLE = 16'h9ffb;
		2602: SAMPLE = 16'h9fd9;
		2603: SAMPLE = 16'h9fb8;
		2604: SAMPLE = 16'h9f97;
		2605: SAMPLE = 16'h9f76;
		2606: SAMPLE = 16'h9f55;
		2607: SAMPLE = 16'h9f34;
		2608: SAMPLE = 16'h9f13;
		2609: SAMPLE = 16'h9ef2;
		2610: SAMPLE = 16'h9ed2;
		2611: SAMPLE = 16'h9eb1;
		2612: SAMPLE = 16'h9e90;
		2613: SAMPLE = 16'h9e70;
		2614: SAMPLE = 16'h9e4f;
		2615: SAMPLE = 16'h9e2f;
		2616: SAMPLE = 16'h9e0e;
		2617: SAMPLE = 16'h9dee;
		2618: SAMPLE = 16'h9dce;
		2619: SAMPLE = 16'h9dae;
		2620: SAMPLE = 16'h9d8e;
		2621: SAMPLE = 16'h9d6d;
		2622: SAMPLE = 16'h9d4d;
		2623: SAMPLE = 16'h9d2d;
		2624: SAMPLE = 16'h9d0d;
		2625: SAMPLE = 16'h9cee;
		2626: SAMPLE = 16'h9cce;
		2627: SAMPLE = 16'h9cae;
		2628: SAMPLE = 16'h9c8e;
		2629: SAMPLE = 16'h9c6f;
		2630: SAMPLE = 16'h9c4f;
		2631: SAMPLE = 16'h9c30;
		2632: SAMPLE = 16'h9c10;
		2633: SAMPLE = 16'h9bf1;
		2634: SAMPLE = 16'h9bd2;
		2635: SAMPLE = 16'h9bb2;
		2636: SAMPLE = 16'h9b93;
		2637: SAMPLE = 16'h9b74;
		2638: SAMPLE = 16'h9b55;
		2639: SAMPLE = 16'h9b36;
		2640: SAMPLE = 16'h9b17;
		2641: SAMPLE = 16'h9af8;
		2642: SAMPLE = 16'h9ad9;
		2643: SAMPLE = 16'h9aba;
		2644: SAMPLE = 16'h9a9c;
		2645: SAMPLE = 16'h9a7d;
		2646: SAMPLE = 16'h9a5f;
		2647: SAMPLE = 16'h9a40;
		2648: SAMPLE = 16'h9a22;
		2649: SAMPLE = 16'h9a03;
		2650: SAMPLE = 16'h99e5;
		2651: SAMPLE = 16'h99c6;
		2652: SAMPLE = 16'h99a8;
		2653: SAMPLE = 16'h998a;
		2654: SAMPLE = 16'h996c;
		2655: SAMPLE = 16'h994e;
		2656: SAMPLE = 16'h9930;
		2657: SAMPLE = 16'h9912;
		2658: SAMPLE = 16'h98f4;
		2659: SAMPLE = 16'h98d6;
		2660: SAMPLE = 16'h98b9;
		2661: SAMPLE = 16'h989b;
		2662: SAMPLE = 16'h987d;
		2663: SAMPLE = 16'h9860;
		2664: SAMPLE = 16'h9842;
		2665: SAMPLE = 16'h9825;
		2666: SAMPLE = 16'h9808;
		2667: SAMPLE = 16'h97ea;
		2668: SAMPLE = 16'h97cd;
		2669: SAMPLE = 16'h97b0;
		2670: SAMPLE = 16'h9793;
		2671: SAMPLE = 16'h9776;
		2672: SAMPLE = 16'h9759;
		2673: SAMPLE = 16'h973c;
		2674: SAMPLE = 16'h971f;
		2675: SAMPLE = 16'h9702;
		2676: SAMPLE = 16'h96e6;
		2677: SAMPLE = 16'h96c9;
		2678: SAMPLE = 16'h96ac;
		2679: SAMPLE = 16'h9690;
		2680: SAMPLE = 16'h9673;
		2681: SAMPLE = 16'h9657;
		2682: SAMPLE = 16'h963b;
		2683: SAMPLE = 16'h961e;
		2684: SAMPLE = 16'h9602;
		2685: SAMPLE = 16'h95e6;
		2686: SAMPLE = 16'h95ca;
		2687: SAMPLE = 16'h95ae;
		2688: SAMPLE = 16'h9592;
		2689: SAMPLE = 16'h9576;
		2690: SAMPLE = 16'h955a;
		2691: SAMPLE = 16'h953e;
		2692: SAMPLE = 16'h9523;
		2693: SAMPLE = 16'h9507;
		2694: SAMPLE = 16'h94ec;
		2695: SAMPLE = 16'h94d0;
		2696: SAMPLE = 16'h94b5;
		2697: SAMPLE = 16'h9499;
		2698: SAMPLE = 16'h947e;
		2699: SAMPLE = 16'h9463;
		2700: SAMPLE = 16'h9447;
		2701: SAMPLE = 16'h942c;
		2702: SAMPLE = 16'h9411;
		2703: SAMPLE = 16'h93f6;
		2704: SAMPLE = 16'h93db;
		2705: SAMPLE = 16'h93c0;
		2706: SAMPLE = 16'h93a6;
		2707: SAMPLE = 16'h938b;
		2708: SAMPLE = 16'h9370;
		2709: SAMPLE = 16'h9356;
		2710: SAMPLE = 16'h933b;
		2711: SAMPLE = 16'h9321;
		2712: SAMPLE = 16'h9306;
		2713: SAMPLE = 16'h92ec;
		2714: SAMPLE = 16'h92d2;
		2715: SAMPLE = 16'h92b7;
		2716: SAMPLE = 16'h929d;
		2717: SAMPLE = 16'h9283;
		2718: SAMPLE = 16'h9269;
		2719: SAMPLE = 16'h924f;
		2720: SAMPLE = 16'h9235;
		2721: SAMPLE = 16'h921c;
		2722: SAMPLE = 16'h9202;
		2723: SAMPLE = 16'h91e8;
		2724: SAMPLE = 16'h91cf;
		2725: SAMPLE = 16'h91b5;
		2726: SAMPLE = 16'h919c;
		2727: SAMPLE = 16'h9182;
		2728: SAMPLE = 16'h9169;
		2729: SAMPLE = 16'h9150;
		2730: SAMPLE = 16'h9136;
		2731: SAMPLE = 16'h911d;
		2732: SAMPLE = 16'h9104;
		2733: SAMPLE = 16'h90eb;
		2734: SAMPLE = 16'h90d2;
		2735: SAMPLE = 16'h90b9;
		2736: SAMPLE = 16'h90a0;
		2737: SAMPLE = 16'h9088;
		2738: SAMPLE = 16'h906f;
		2739: SAMPLE = 16'h9056;
		2740: SAMPLE = 16'h903e;
		2741: SAMPLE = 16'h9025;
		2742: SAMPLE = 16'h900d;
		2743: SAMPLE = 16'h8ff5;
		2744: SAMPLE = 16'h8fdc;
		2745: SAMPLE = 16'h8fc4;
		2746: SAMPLE = 16'h8fac;
		2747: SAMPLE = 16'h8f94;
		2748: SAMPLE = 16'h8f7c;
		2749: SAMPLE = 16'h8f64;
		2750: SAMPLE = 16'h8f4c;
		2751: SAMPLE = 16'h8f34;
		2752: SAMPLE = 16'h8f1d;
		2753: SAMPLE = 16'h8f05;
		2754: SAMPLE = 16'h8eed;
		2755: SAMPLE = 16'h8ed6;
		2756: SAMPLE = 16'h8ebe;
		2757: SAMPLE = 16'h8ea7;
		2758: SAMPLE = 16'h8e90;
		2759: SAMPLE = 16'h8e79;
		2760: SAMPLE = 16'h8e61;
		2761: SAMPLE = 16'h8e4a;
		2762: SAMPLE = 16'h8e33;
		2763: SAMPLE = 16'h8e1c;
		2764: SAMPLE = 16'h8e05;
		2765: SAMPLE = 16'h8dee;
		2766: SAMPLE = 16'h8dd8;
		2767: SAMPLE = 16'h8dc1;
		2768: SAMPLE = 16'h8daa;
		2769: SAMPLE = 16'h8d94;
		2770: SAMPLE = 16'h8d7d;
		2771: SAMPLE = 16'h8d67;
		2772: SAMPLE = 16'h8d50;
		2773: SAMPLE = 16'h8d3a;
		2774: SAMPLE = 16'h8d24;
		2775: SAMPLE = 16'h8d0e;
		2776: SAMPLE = 16'h8cf8;
		2777: SAMPLE = 16'h8ce2;
		2778: SAMPLE = 16'h8ccc;
		2779: SAMPLE = 16'h8cb6;
		2780: SAMPLE = 16'h8ca0;
		2781: SAMPLE = 16'h8c8a;
		2782: SAMPLE = 16'h8c75;
		2783: SAMPLE = 16'h8c5f;
		2784: SAMPLE = 16'h8c4a;
		2785: SAMPLE = 16'h8c34;
		2786: SAMPLE = 16'h8c1f;
		2787: SAMPLE = 16'h8c09;
		2788: SAMPLE = 16'h8bf4;
		2789: SAMPLE = 16'h8bdf;
		2790: SAMPLE = 16'h8bca;
		2791: SAMPLE = 16'h8bb5;
		2792: SAMPLE = 16'h8ba0;
		2793: SAMPLE = 16'h8b8b;
		2794: SAMPLE = 16'h8b76;
		2795: SAMPLE = 16'h8b61;
		2796: SAMPLE = 16'h8b4d;
		2797: SAMPLE = 16'h8b38;
		2798: SAMPLE = 16'h8b24;
		2799: SAMPLE = 16'h8b0f;
		2800: SAMPLE = 16'h8afb;
		2801: SAMPLE = 16'h8ae6;
		2802: SAMPLE = 16'h8ad2;
		2803: SAMPLE = 16'h8abe;
		2804: SAMPLE = 16'h8aaa;
		2805: SAMPLE = 16'h8a96;
		2806: SAMPLE = 16'h8a82;
		2807: SAMPLE = 16'h8a6e;
		2808: SAMPLE = 16'h8a5a;
		2809: SAMPLE = 16'h8a46;
		2810: SAMPLE = 16'h8a33;
		2811: SAMPLE = 16'h8a1f;
		2812: SAMPLE = 16'h8a0b;
		2813: SAMPLE = 16'h89f8;
		2814: SAMPLE = 16'h89e4;
		2815: SAMPLE = 16'h89d1;
		2816: SAMPLE = 16'h89be;
		2817: SAMPLE = 16'h89ab;
		2818: SAMPLE = 16'h8997;
		2819: SAMPLE = 16'h8984;
		2820: SAMPLE = 16'h8971;
		2821: SAMPLE = 16'h895f;
		2822: SAMPLE = 16'h894c;
		2823: SAMPLE = 16'h8939;
		2824: SAMPLE = 16'h8926;
		2825: SAMPLE = 16'h8914;
		2826: SAMPLE = 16'h8901;
		2827: SAMPLE = 16'h88ef;
		2828: SAMPLE = 16'h88dc;
		2829: SAMPLE = 16'h88ca;
		2830: SAMPLE = 16'h88b8;
		2831: SAMPLE = 16'h88a5;
		2832: SAMPLE = 16'h8893;
		2833: SAMPLE = 16'h8881;
		2834: SAMPLE = 16'h886f;
		2835: SAMPLE = 16'h885d;
		2836: SAMPLE = 16'h884b;
		2837: SAMPLE = 16'h883a;
		2838: SAMPLE = 16'h8828;
		2839: SAMPLE = 16'h8816;
		2840: SAMPLE = 16'h8805;
		2841: SAMPLE = 16'h87f3;
		2842: SAMPLE = 16'h87e2;
		2843: SAMPLE = 16'h87d1;
		2844: SAMPLE = 16'h87bf;
		2845: SAMPLE = 16'h87ae;
		2846: SAMPLE = 16'h879d;
		2847: SAMPLE = 16'h878c;
		2848: SAMPLE = 16'h877b;
		2849: SAMPLE = 16'h876a;
		2850: SAMPLE = 16'h8759;
		2851: SAMPLE = 16'h8749;
		2852: SAMPLE = 16'h8738;
		2853: SAMPLE = 16'h8727;
		2854: SAMPLE = 16'h8717;
		2855: SAMPLE = 16'h8706;
		2856: SAMPLE = 16'h86f6;
		2857: SAMPLE = 16'h86e6;
		2858: SAMPLE = 16'h86d5;
		2859: SAMPLE = 16'h86c5;
		2860: SAMPLE = 16'h86b5;
		2861: SAMPLE = 16'h86a5;
		2862: SAMPLE = 16'h8695;
		2863: SAMPLE = 16'h8685;
		2864: SAMPLE = 16'h8675;
		2865: SAMPLE = 16'h8666;
		2866: SAMPLE = 16'h8656;
		2867: SAMPLE = 16'h8646;
		2868: SAMPLE = 16'h8637;
		2869: SAMPLE = 16'h8627;
		2870: SAMPLE = 16'h8618;
		2871: SAMPLE = 16'h8609;
		2872: SAMPLE = 16'h85fa;
		2873: SAMPLE = 16'h85ea;
		2874: SAMPLE = 16'h85db;
		2875: SAMPLE = 16'h85cc;
		2876: SAMPLE = 16'h85bd;
		2877: SAMPLE = 16'h85af;
		2878: SAMPLE = 16'h85a0;
		2879: SAMPLE = 16'h8591;
		2880: SAMPLE = 16'h8582;
		2881: SAMPLE = 16'h8574;
		2882: SAMPLE = 16'h8565;
		2883: SAMPLE = 16'h8557;
		2884: SAMPLE = 16'h8549;
		2885: SAMPLE = 16'h853a;
		2886: SAMPLE = 16'h852c;
		2887: SAMPLE = 16'h851e;
		2888: SAMPLE = 16'h8510;
		2889: SAMPLE = 16'h8502;
		2890: SAMPLE = 16'h84f4;
		2891: SAMPLE = 16'h84e6;
		2892: SAMPLE = 16'h84d9;
		2893: SAMPLE = 16'h84cb;
		2894: SAMPLE = 16'h84bd;
		2895: SAMPLE = 16'h84b0;
		2896: SAMPLE = 16'h84a2;
		2897: SAMPLE = 16'h8495;
		2898: SAMPLE = 16'h8488;
		2899: SAMPLE = 16'h847b;
		2900: SAMPLE = 16'h846d;
		2901: SAMPLE = 16'h8460;
		2902: SAMPLE = 16'h8453;
		2903: SAMPLE = 16'h8446;
		2904: SAMPLE = 16'h843a;
		2905: SAMPLE = 16'h842d;
		2906: SAMPLE = 16'h8420;
		2907: SAMPLE = 16'h8414;
		2908: SAMPLE = 16'h8407;
		2909: SAMPLE = 16'h83fa;
		2910: SAMPLE = 16'h83ee;
		2911: SAMPLE = 16'h83e2;
		2912: SAMPLE = 16'h83d6;
		2913: SAMPLE = 16'h83c9;
		2914: SAMPLE = 16'h83bd;
		2915: SAMPLE = 16'h83b1;
		2916: SAMPLE = 16'h83a5;
		2917: SAMPLE = 16'h8399;
		2918: SAMPLE = 16'h838e;
		2919: SAMPLE = 16'h8382;
		2920: SAMPLE = 16'h8376;
		2921: SAMPLE = 16'h836b;
		2922: SAMPLE = 16'h835f;
		2923: SAMPLE = 16'h8354;
		2924: SAMPLE = 16'h8348;
		2925: SAMPLE = 16'h833d;
		2926: SAMPLE = 16'h8332;
		2927: SAMPLE = 16'h8327;
		2928: SAMPLE = 16'h831c;
		2929: SAMPLE = 16'h8311;
		2930: SAMPLE = 16'h8306;
		2931: SAMPLE = 16'h82fb;
		2932: SAMPLE = 16'h82f0;
		2933: SAMPLE = 16'h82e6;
		2934: SAMPLE = 16'h82db;
		2935: SAMPLE = 16'h82d0;
		2936: SAMPLE = 16'h82c6;
		2937: SAMPLE = 16'h82bc;
		2938: SAMPLE = 16'h82b1;
		2939: SAMPLE = 16'h82a7;
		2940: SAMPLE = 16'h829d;
		2941: SAMPLE = 16'h8293;
		2942: SAMPLE = 16'h8289;
		2943: SAMPLE = 16'h827f;
		2944: SAMPLE = 16'h8275;
		2945: SAMPLE = 16'h826b;
		2946: SAMPLE = 16'h8262;
		2947: SAMPLE = 16'h8258;
		2948: SAMPLE = 16'h824f;
		2949: SAMPLE = 16'h8245;
		2950: SAMPLE = 16'h823c;
		2951: SAMPLE = 16'h8232;
		2952: SAMPLE = 16'h8229;
		2953: SAMPLE = 16'h8220;
		2954: SAMPLE = 16'h8217;
		2955: SAMPLE = 16'h820e;
		2956: SAMPLE = 16'h8205;
		2957: SAMPLE = 16'h81fc;
		2958: SAMPLE = 16'h81f3;
		2959: SAMPLE = 16'h81eb;
		2960: SAMPLE = 16'h81e2;
		2961: SAMPLE = 16'h81d9;
		2962: SAMPLE = 16'h81d1;
		2963: SAMPLE = 16'h81c8;
		2964: SAMPLE = 16'h81c0;
		2965: SAMPLE = 16'h81b8;
		2966: SAMPLE = 16'h81b0;
		2967: SAMPLE = 16'h81a8;
		2968: SAMPLE = 16'h81a0;
		2969: SAMPLE = 16'h8198;
		2970: SAMPLE = 16'h8190;
		2971: SAMPLE = 16'h8188;
		2972: SAMPLE = 16'h8180;
		2973: SAMPLE = 16'h8179;
		2974: SAMPLE = 16'h8171;
		2975: SAMPLE = 16'h816a;
		2976: SAMPLE = 16'h8162;
		2977: SAMPLE = 16'h815b;
		2978: SAMPLE = 16'h8154;
		2979: SAMPLE = 16'h814c;
		2980: SAMPLE = 16'h8145;
		2981: SAMPLE = 16'h813e;
		2982: SAMPLE = 16'h8137;
		2983: SAMPLE = 16'h8130;
		2984: SAMPLE = 16'h812a;
		2985: SAMPLE = 16'h8123;
		2986: SAMPLE = 16'h811c;
		2987: SAMPLE = 16'h8116;
		2988: SAMPLE = 16'h810f;
		2989: SAMPLE = 16'h8109;
		2990: SAMPLE = 16'h8102;
		2991: SAMPLE = 16'h80fc;
		2992: SAMPLE = 16'h80f6;
		2993: SAMPLE = 16'h80f0;
		2994: SAMPLE = 16'h80ea;
		2995: SAMPLE = 16'h80e4;
		2996: SAMPLE = 16'h80de;
		2997: SAMPLE = 16'h80d8;
		2998: SAMPLE = 16'h80d2;
		2999: SAMPLE = 16'h80cd;
		3000: SAMPLE = 16'h80c7;
		3001: SAMPLE = 16'h80c2;
		3002: SAMPLE = 16'h80bc;
		3003: SAMPLE = 16'h80b7;
		3004: SAMPLE = 16'h80b2;
		3005: SAMPLE = 16'h80ac;
		3006: SAMPLE = 16'h80a7;
		3007: SAMPLE = 16'h80a2;
		3008: SAMPLE = 16'h809d;
		3009: SAMPLE = 16'h8098;
		3010: SAMPLE = 16'h8094;
		3011: SAMPLE = 16'h808f;
		3012: SAMPLE = 16'h808a;
		3013: SAMPLE = 16'h8086;
		3014: SAMPLE = 16'h8081;
		3015: SAMPLE = 16'h807d;
		3016: SAMPLE = 16'h8078;
		3017: SAMPLE = 16'h8074;
		3018: SAMPLE = 16'h8070;
		3019: SAMPLE = 16'h806c;
		3020: SAMPLE = 16'h8068;
		3021: SAMPLE = 16'h8064;
		3022: SAMPLE = 16'h8060;
		3023: SAMPLE = 16'h805c;
		3024: SAMPLE = 16'h8058;
		3025: SAMPLE = 16'h8055;
		3026: SAMPLE = 16'h8051;
		3027: SAMPLE = 16'h804e;
		3028: SAMPLE = 16'h804a;
		3029: SAMPLE = 16'h8047;
		3030: SAMPLE = 16'h8043;
		3031: SAMPLE = 16'h8040;
		3032: SAMPLE = 16'h803d;
		3033: SAMPLE = 16'h803a;
		3034: SAMPLE = 16'h8037;
		3035: SAMPLE = 16'h8034;
		3036: SAMPLE = 16'h8031;
		3037: SAMPLE = 16'h802f;
		3038: SAMPLE = 16'h802c;
		3039: SAMPLE = 16'h8029;
		3040: SAMPLE = 16'h8027;
		3041: SAMPLE = 16'h8025;
		3042: SAMPLE = 16'h8022;
		3043: SAMPLE = 16'h8020;
		3044: SAMPLE = 16'h801e;
		3045: SAMPLE = 16'h801c;
		3046: SAMPLE = 16'h801a;
		3047: SAMPLE = 16'h8018;
		3048: SAMPLE = 16'h8016;
		3049: SAMPLE = 16'h8014;
		3050: SAMPLE = 16'h8012;
		3051: SAMPLE = 16'h8011;
		3052: SAMPLE = 16'h800f;
		3053: SAMPLE = 16'h800d;
		3054: SAMPLE = 16'h800c;
		3055: SAMPLE = 16'h800b;
		3056: SAMPLE = 16'h8009;
		3057: SAMPLE = 16'h8008;
		3058: SAMPLE = 16'h8007;
		3059: SAMPLE = 16'h8006;
		3060: SAMPLE = 16'h8005;
		3061: SAMPLE = 16'h8004;
		3062: SAMPLE = 16'h8003;
		3063: SAMPLE = 16'h8003;
		3064: SAMPLE = 16'h8002;
		3065: SAMPLE = 16'h8001;
		3066: SAMPLE = 16'h8001;
		3067: SAMPLE = 16'h8000;
		3068: SAMPLE = 16'h8000;
		3069: SAMPLE = 16'h8000;
		3070: SAMPLE = 16'h8000;
		3071: SAMPLE = 16'h8000;
		3072: SAMPLE = 16'h8000;
		3073: SAMPLE = 16'h8000;
		3074: SAMPLE = 16'h8000;
		3075: SAMPLE = 16'h8000;
		3076: SAMPLE = 16'h8000;
		3077: SAMPLE = 16'h8000;
		3078: SAMPLE = 16'h8001;
		3079: SAMPLE = 16'h8001;
		3080: SAMPLE = 16'h8002;
		3081: SAMPLE = 16'h8003;
		3082: SAMPLE = 16'h8003;
		3083: SAMPLE = 16'h8004;
		3084: SAMPLE = 16'h8005;
		3085: SAMPLE = 16'h8006;
		3086: SAMPLE = 16'h8007;
		3087: SAMPLE = 16'h8008;
		3088: SAMPLE = 16'h8009;
		3089: SAMPLE = 16'h800b;
		3090: SAMPLE = 16'h800c;
		3091: SAMPLE = 16'h800d;
		3092: SAMPLE = 16'h800f;
		3093: SAMPLE = 16'h8011;
		3094: SAMPLE = 16'h8012;
		3095: SAMPLE = 16'h8014;
		3096: SAMPLE = 16'h8016;
		3097: SAMPLE = 16'h8018;
		3098: SAMPLE = 16'h801a;
		3099: SAMPLE = 16'h801c;
		3100: SAMPLE = 16'h801e;
		3101: SAMPLE = 16'h8020;
		3102: SAMPLE = 16'h8022;
		3103: SAMPLE = 16'h8025;
		3104: SAMPLE = 16'h8027;
		3105: SAMPLE = 16'h8029;
		3106: SAMPLE = 16'h802c;
		3107: SAMPLE = 16'h802f;
		3108: SAMPLE = 16'h8031;
		3109: SAMPLE = 16'h8034;
		3110: SAMPLE = 16'h8037;
		3111: SAMPLE = 16'h803a;
		3112: SAMPLE = 16'h803d;
		3113: SAMPLE = 16'h8040;
		3114: SAMPLE = 16'h8043;
		3115: SAMPLE = 16'h8047;
		3116: SAMPLE = 16'h804a;
		3117: SAMPLE = 16'h804e;
		3118: SAMPLE = 16'h8051;
		3119: SAMPLE = 16'h8055;
		3120: SAMPLE = 16'h8058;
		3121: SAMPLE = 16'h805c;
		3122: SAMPLE = 16'h8060;
		3123: SAMPLE = 16'h8064;
		3124: SAMPLE = 16'h8068;
		3125: SAMPLE = 16'h806c;
		3126: SAMPLE = 16'h8070;
		3127: SAMPLE = 16'h8074;
		3128: SAMPLE = 16'h8078;
		3129: SAMPLE = 16'h807d;
		3130: SAMPLE = 16'h8081;
		3131: SAMPLE = 16'h8086;
		3132: SAMPLE = 16'h808a;
		3133: SAMPLE = 16'h808f;
		3134: SAMPLE = 16'h8094;
		3135: SAMPLE = 16'h8098;
		3136: SAMPLE = 16'h809d;
		3137: SAMPLE = 16'h80a2;
		3138: SAMPLE = 16'h80a7;
		3139: SAMPLE = 16'h80ac;
		3140: SAMPLE = 16'h80b2;
		3141: SAMPLE = 16'h80b7;
		3142: SAMPLE = 16'h80bc;
		3143: SAMPLE = 16'h80c2;
		3144: SAMPLE = 16'h80c7;
		3145: SAMPLE = 16'h80cd;
		3146: SAMPLE = 16'h80d2;
		3147: SAMPLE = 16'h80d8;
		3148: SAMPLE = 16'h80de;
		3149: SAMPLE = 16'h80e4;
		3150: SAMPLE = 16'h80ea;
		3151: SAMPLE = 16'h80f0;
		3152: SAMPLE = 16'h80f6;
		3153: SAMPLE = 16'h80fc;
		3154: SAMPLE = 16'h8102;
		3155: SAMPLE = 16'h8109;
		3156: SAMPLE = 16'h810f;
		3157: SAMPLE = 16'h8116;
		3158: SAMPLE = 16'h811c;
		3159: SAMPLE = 16'h8123;
		3160: SAMPLE = 16'h812a;
		3161: SAMPLE = 16'h8130;
		3162: SAMPLE = 16'h8137;
		3163: SAMPLE = 16'h813e;
		3164: SAMPLE = 16'h8145;
		3165: SAMPLE = 16'h814c;
		3166: SAMPLE = 16'h8154;
		3167: SAMPLE = 16'h815b;
		3168: SAMPLE = 16'h8162;
		3169: SAMPLE = 16'h816a;
		3170: SAMPLE = 16'h8171;
		3171: SAMPLE = 16'h8179;
		3172: SAMPLE = 16'h8180;
		3173: SAMPLE = 16'h8188;
		3174: SAMPLE = 16'h8190;
		3175: SAMPLE = 16'h8198;
		3176: SAMPLE = 16'h81a0;
		3177: SAMPLE = 16'h81a8;
		3178: SAMPLE = 16'h81b0;
		3179: SAMPLE = 16'h81b8;
		3180: SAMPLE = 16'h81c0;
		3181: SAMPLE = 16'h81c8;
		3182: SAMPLE = 16'h81d1;
		3183: SAMPLE = 16'h81d9;
		3184: SAMPLE = 16'h81e2;
		3185: SAMPLE = 16'h81eb;
		3186: SAMPLE = 16'h81f3;
		3187: SAMPLE = 16'h81fc;
		3188: SAMPLE = 16'h8205;
		3189: SAMPLE = 16'h820e;
		3190: SAMPLE = 16'h8217;
		3191: SAMPLE = 16'h8220;
		3192: SAMPLE = 16'h8229;
		3193: SAMPLE = 16'h8232;
		3194: SAMPLE = 16'h823c;
		3195: SAMPLE = 16'h8245;
		3196: SAMPLE = 16'h824f;
		3197: SAMPLE = 16'h8258;
		3198: SAMPLE = 16'h8262;
		3199: SAMPLE = 16'h826b;
		3200: SAMPLE = 16'h8275;
		3201: SAMPLE = 16'h827f;
		3202: SAMPLE = 16'h8289;
		3203: SAMPLE = 16'h8293;
		3204: SAMPLE = 16'h829d;
		3205: SAMPLE = 16'h82a7;
		3206: SAMPLE = 16'h82b1;
		3207: SAMPLE = 16'h82bc;
		3208: SAMPLE = 16'h82c6;
		3209: SAMPLE = 16'h82d0;
		3210: SAMPLE = 16'h82db;
		3211: SAMPLE = 16'h82e6;
		3212: SAMPLE = 16'h82f0;
		3213: SAMPLE = 16'h82fb;
		3214: SAMPLE = 16'h8306;
		3215: SAMPLE = 16'h8311;
		3216: SAMPLE = 16'h831c;
		3217: SAMPLE = 16'h8327;
		3218: SAMPLE = 16'h8332;
		3219: SAMPLE = 16'h833d;
		3220: SAMPLE = 16'h8348;
		3221: SAMPLE = 16'h8354;
		3222: SAMPLE = 16'h835f;
		3223: SAMPLE = 16'h836b;
		3224: SAMPLE = 16'h8376;
		3225: SAMPLE = 16'h8382;
		3226: SAMPLE = 16'h838e;
		3227: SAMPLE = 16'h8399;
		3228: SAMPLE = 16'h83a5;
		3229: SAMPLE = 16'h83b1;
		3230: SAMPLE = 16'h83bd;
		3231: SAMPLE = 16'h83c9;
		3232: SAMPLE = 16'h83d6;
		3233: SAMPLE = 16'h83e2;
		3234: SAMPLE = 16'h83ee;
		3235: SAMPLE = 16'h83fa;
		3236: SAMPLE = 16'h8407;
		3237: SAMPLE = 16'h8414;
		3238: SAMPLE = 16'h8420;
		3239: SAMPLE = 16'h842d;
		3240: SAMPLE = 16'h843a;
		3241: SAMPLE = 16'h8446;
		3242: SAMPLE = 16'h8453;
		3243: SAMPLE = 16'h8460;
		3244: SAMPLE = 16'h846d;
		3245: SAMPLE = 16'h847b;
		3246: SAMPLE = 16'h8488;
		3247: SAMPLE = 16'h8495;
		3248: SAMPLE = 16'h84a2;
		3249: SAMPLE = 16'h84b0;
		3250: SAMPLE = 16'h84bd;
		3251: SAMPLE = 16'h84cb;
		3252: SAMPLE = 16'h84d9;
		3253: SAMPLE = 16'h84e6;
		3254: SAMPLE = 16'h84f4;
		3255: SAMPLE = 16'h8502;
		3256: SAMPLE = 16'h8510;
		3257: SAMPLE = 16'h851e;
		3258: SAMPLE = 16'h852c;
		3259: SAMPLE = 16'h853a;
		3260: SAMPLE = 16'h8549;
		3261: SAMPLE = 16'h8557;
		3262: SAMPLE = 16'h8565;
		3263: SAMPLE = 16'h8574;
		3264: SAMPLE = 16'h8582;
		3265: SAMPLE = 16'h8591;
		3266: SAMPLE = 16'h85a0;
		3267: SAMPLE = 16'h85af;
		3268: SAMPLE = 16'h85bd;
		3269: SAMPLE = 16'h85cc;
		3270: SAMPLE = 16'h85db;
		3271: SAMPLE = 16'h85ea;
		3272: SAMPLE = 16'h85fa;
		3273: SAMPLE = 16'h8609;
		3274: SAMPLE = 16'h8618;
		3275: SAMPLE = 16'h8627;
		3276: SAMPLE = 16'h8637;
		3277: SAMPLE = 16'h8646;
		3278: SAMPLE = 16'h8656;
		3279: SAMPLE = 16'h8666;
		3280: SAMPLE = 16'h8675;
		3281: SAMPLE = 16'h8685;
		3282: SAMPLE = 16'h8695;
		3283: SAMPLE = 16'h86a5;
		3284: SAMPLE = 16'h86b5;
		3285: SAMPLE = 16'h86c5;
		3286: SAMPLE = 16'h86d5;
		3287: SAMPLE = 16'h86e6;
		3288: SAMPLE = 16'h86f6;
		3289: SAMPLE = 16'h8706;
		3290: SAMPLE = 16'h8717;
		3291: SAMPLE = 16'h8727;
		3292: SAMPLE = 16'h8738;
		3293: SAMPLE = 16'h8749;
		3294: SAMPLE = 16'h8759;
		3295: SAMPLE = 16'h876a;
		3296: SAMPLE = 16'h877b;
		3297: SAMPLE = 16'h878c;
		3298: SAMPLE = 16'h879d;
		3299: SAMPLE = 16'h87ae;
		3300: SAMPLE = 16'h87bf;
		3301: SAMPLE = 16'h87d1;
		3302: SAMPLE = 16'h87e2;
		3303: SAMPLE = 16'h87f3;
		3304: SAMPLE = 16'h8805;
		3305: SAMPLE = 16'h8816;
		3306: SAMPLE = 16'h8828;
		3307: SAMPLE = 16'h883a;
		3308: SAMPLE = 16'h884b;
		3309: SAMPLE = 16'h885d;
		3310: SAMPLE = 16'h886f;
		3311: SAMPLE = 16'h8881;
		3312: SAMPLE = 16'h8893;
		3313: SAMPLE = 16'h88a5;
		3314: SAMPLE = 16'h88b8;
		3315: SAMPLE = 16'h88ca;
		3316: SAMPLE = 16'h88dc;
		3317: SAMPLE = 16'h88ef;
		3318: SAMPLE = 16'h8901;
		3319: SAMPLE = 16'h8914;
		3320: SAMPLE = 16'h8926;
		3321: SAMPLE = 16'h8939;
		3322: SAMPLE = 16'h894c;
		3323: SAMPLE = 16'h895f;
		3324: SAMPLE = 16'h8971;
		3325: SAMPLE = 16'h8984;
		3326: SAMPLE = 16'h8997;
		3327: SAMPLE = 16'h89ab;
		3328: SAMPLE = 16'h89be;
		3329: SAMPLE = 16'h89d1;
		3330: SAMPLE = 16'h89e4;
		3331: SAMPLE = 16'h89f8;
		3332: SAMPLE = 16'h8a0b;
		3333: SAMPLE = 16'h8a1f;
		3334: SAMPLE = 16'h8a33;
		3335: SAMPLE = 16'h8a46;
		3336: SAMPLE = 16'h8a5a;
		3337: SAMPLE = 16'h8a6e;
		3338: SAMPLE = 16'h8a82;
		3339: SAMPLE = 16'h8a96;
		3340: SAMPLE = 16'h8aaa;
		3341: SAMPLE = 16'h8abe;
		3342: SAMPLE = 16'h8ad2;
		3343: SAMPLE = 16'h8ae6;
		3344: SAMPLE = 16'h8afb;
		3345: SAMPLE = 16'h8b0f;
		3346: SAMPLE = 16'h8b24;
		3347: SAMPLE = 16'h8b38;
		3348: SAMPLE = 16'h8b4d;
		3349: SAMPLE = 16'h8b61;
		3350: SAMPLE = 16'h8b76;
		3351: SAMPLE = 16'h8b8b;
		3352: SAMPLE = 16'h8ba0;
		3353: SAMPLE = 16'h8bb5;
		3354: SAMPLE = 16'h8bca;
		3355: SAMPLE = 16'h8bdf;
		3356: SAMPLE = 16'h8bf4;
		3357: SAMPLE = 16'h8c09;
		3358: SAMPLE = 16'h8c1f;
		3359: SAMPLE = 16'h8c34;
		3360: SAMPLE = 16'h8c4a;
		3361: SAMPLE = 16'h8c5f;
		3362: SAMPLE = 16'h8c75;
		3363: SAMPLE = 16'h8c8a;
		3364: SAMPLE = 16'h8ca0;
		3365: SAMPLE = 16'h8cb6;
		3366: SAMPLE = 16'h8ccc;
		3367: SAMPLE = 16'h8ce2;
		3368: SAMPLE = 16'h8cf8;
		3369: SAMPLE = 16'h8d0e;
		3370: SAMPLE = 16'h8d24;
		3371: SAMPLE = 16'h8d3a;
		3372: SAMPLE = 16'h8d50;
		3373: SAMPLE = 16'h8d67;
		3374: SAMPLE = 16'h8d7d;
		3375: SAMPLE = 16'h8d94;
		3376: SAMPLE = 16'h8daa;
		3377: SAMPLE = 16'h8dc1;
		3378: SAMPLE = 16'h8dd8;
		3379: SAMPLE = 16'h8dee;
		3380: SAMPLE = 16'h8e05;
		3381: SAMPLE = 16'h8e1c;
		3382: SAMPLE = 16'h8e33;
		3383: SAMPLE = 16'h8e4a;
		3384: SAMPLE = 16'h8e61;
		3385: SAMPLE = 16'h8e79;
		3386: SAMPLE = 16'h8e90;
		3387: SAMPLE = 16'h8ea7;
		3388: SAMPLE = 16'h8ebe;
		3389: SAMPLE = 16'h8ed6;
		3390: SAMPLE = 16'h8eed;
		3391: SAMPLE = 16'h8f05;
		3392: SAMPLE = 16'h8f1d;
		3393: SAMPLE = 16'h8f34;
		3394: SAMPLE = 16'h8f4c;
		3395: SAMPLE = 16'h8f64;
		3396: SAMPLE = 16'h8f7c;
		3397: SAMPLE = 16'h8f94;
		3398: SAMPLE = 16'h8fac;
		3399: SAMPLE = 16'h8fc4;
		3400: SAMPLE = 16'h8fdc;
		3401: SAMPLE = 16'h8ff5;
		3402: SAMPLE = 16'h900d;
		3403: SAMPLE = 16'h9025;
		3404: SAMPLE = 16'h903e;
		3405: SAMPLE = 16'h9056;
		3406: SAMPLE = 16'h906f;
		3407: SAMPLE = 16'h9088;
		3408: SAMPLE = 16'h90a0;
		3409: SAMPLE = 16'h90b9;
		3410: SAMPLE = 16'h90d2;
		3411: SAMPLE = 16'h90eb;
		3412: SAMPLE = 16'h9104;
		3413: SAMPLE = 16'h911d;
		3414: SAMPLE = 16'h9136;
		3415: SAMPLE = 16'h9150;
		3416: SAMPLE = 16'h9169;
		3417: SAMPLE = 16'h9182;
		3418: SAMPLE = 16'h919c;
		3419: SAMPLE = 16'h91b5;
		3420: SAMPLE = 16'h91cf;
		3421: SAMPLE = 16'h91e8;
		3422: SAMPLE = 16'h9202;
		3423: SAMPLE = 16'h921c;
		3424: SAMPLE = 16'h9235;
		3425: SAMPLE = 16'h924f;
		3426: SAMPLE = 16'h9269;
		3427: SAMPLE = 16'h9283;
		3428: SAMPLE = 16'h929d;
		3429: SAMPLE = 16'h92b7;
		3430: SAMPLE = 16'h92d2;
		3431: SAMPLE = 16'h92ec;
		3432: SAMPLE = 16'h9306;
		3433: SAMPLE = 16'h9321;
		3434: SAMPLE = 16'h933b;
		3435: SAMPLE = 16'h9356;
		3436: SAMPLE = 16'h9370;
		3437: SAMPLE = 16'h938b;
		3438: SAMPLE = 16'h93a6;
		3439: SAMPLE = 16'h93c0;
		3440: SAMPLE = 16'h93db;
		3441: SAMPLE = 16'h93f6;
		3442: SAMPLE = 16'h9411;
		3443: SAMPLE = 16'h942c;
		3444: SAMPLE = 16'h9447;
		3445: SAMPLE = 16'h9463;
		3446: SAMPLE = 16'h947e;
		3447: SAMPLE = 16'h9499;
		3448: SAMPLE = 16'h94b5;
		3449: SAMPLE = 16'h94d0;
		3450: SAMPLE = 16'h94ec;
		3451: SAMPLE = 16'h9507;
		3452: SAMPLE = 16'h9523;
		3453: SAMPLE = 16'h953e;
		3454: SAMPLE = 16'h955a;
		3455: SAMPLE = 16'h9576;
		3456: SAMPLE = 16'h9592;
		3457: SAMPLE = 16'h95ae;
		3458: SAMPLE = 16'h95ca;
		3459: SAMPLE = 16'h95e6;
		3460: SAMPLE = 16'h9602;
		3461: SAMPLE = 16'h961e;
		3462: SAMPLE = 16'h963b;
		3463: SAMPLE = 16'h9657;
		3464: SAMPLE = 16'h9673;
		3465: SAMPLE = 16'h9690;
		3466: SAMPLE = 16'h96ac;
		3467: SAMPLE = 16'h96c9;
		3468: SAMPLE = 16'h96e6;
		3469: SAMPLE = 16'h9702;
		3470: SAMPLE = 16'h971f;
		3471: SAMPLE = 16'h973c;
		3472: SAMPLE = 16'h9759;
		3473: SAMPLE = 16'h9776;
		3474: SAMPLE = 16'h9793;
		3475: SAMPLE = 16'h97b0;
		3476: SAMPLE = 16'h97cd;
		3477: SAMPLE = 16'h97ea;
		3478: SAMPLE = 16'h9808;
		3479: SAMPLE = 16'h9825;
		3480: SAMPLE = 16'h9842;
		3481: SAMPLE = 16'h9860;
		3482: SAMPLE = 16'h987d;
		3483: SAMPLE = 16'h989b;
		3484: SAMPLE = 16'h98b9;
		3485: SAMPLE = 16'h98d6;
		3486: SAMPLE = 16'h98f4;
		3487: SAMPLE = 16'h9912;
		3488: SAMPLE = 16'h9930;
		3489: SAMPLE = 16'h994e;
		3490: SAMPLE = 16'h996c;
		3491: SAMPLE = 16'h998a;
		3492: SAMPLE = 16'h99a8;
		3493: SAMPLE = 16'h99c6;
		3494: SAMPLE = 16'h99e5;
		3495: SAMPLE = 16'h9a03;
		3496: SAMPLE = 16'h9a22;
		3497: SAMPLE = 16'h9a40;
		3498: SAMPLE = 16'h9a5f;
		3499: SAMPLE = 16'h9a7d;
		3500: SAMPLE = 16'h9a9c;
		3501: SAMPLE = 16'h9aba;
		3502: SAMPLE = 16'h9ad9;
		3503: SAMPLE = 16'h9af8;
		3504: SAMPLE = 16'h9b17;
		3505: SAMPLE = 16'h9b36;
		3506: SAMPLE = 16'h9b55;
		3507: SAMPLE = 16'h9b74;
		3508: SAMPLE = 16'h9b93;
		3509: SAMPLE = 16'h9bb2;
		3510: SAMPLE = 16'h9bd2;
		3511: SAMPLE = 16'h9bf1;
		3512: SAMPLE = 16'h9c10;
		3513: SAMPLE = 16'h9c30;
		3514: SAMPLE = 16'h9c4f;
		3515: SAMPLE = 16'h9c6f;
		3516: SAMPLE = 16'h9c8e;
		3517: SAMPLE = 16'h9cae;
		3518: SAMPLE = 16'h9cce;
		3519: SAMPLE = 16'h9cee;
		3520: SAMPLE = 16'h9d0d;
		3521: SAMPLE = 16'h9d2d;
		3522: SAMPLE = 16'h9d4d;
		3523: SAMPLE = 16'h9d6d;
		3524: SAMPLE = 16'h9d8e;
		3525: SAMPLE = 16'h9dae;
		3526: SAMPLE = 16'h9dce;
		3527: SAMPLE = 16'h9dee;
		3528: SAMPLE = 16'h9e0e;
		3529: SAMPLE = 16'h9e2f;
		3530: SAMPLE = 16'h9e4f;
		3531: SAMPLE = 16'h9e70;
		3532: SAMPLE = 16'h9e90;
		3533: SAMPLE = 16'h9eb1;
		3534: SAMPLE = 16'h9ed2;
		3535: SAMPLE = 16'h9ef2;
		3536: SAMPLE = 16'h9f13;
		3537: SAMPLE = 16'h9f34;
		3538: SAMPLE = 16'h9f55;
		3539: SAMPLE = 16'h9f76;
		3540: SAMPLE = 16'h9f97;
		3541: SAMPLE = 16'h9fb8;
		3542: SAMPLE = 16'h9fd9;
		3543: SAMPLE = 16'h9ffb;
		3544: SAMPLE = 16'ha01c;
		3545: SAMPLE = 16'ha03d;
		3546: SAMPLE = 16'ha05f;
		3547: SAMPLE = 16'ha080;
		3548: SAMPLE = 16'ha0a1;
		3549: SAMPLE = 16'ha0c3;
		3550: SAMPLE = 16'ha0e5;
		3551: SAMPLE = 16'ha106;
		3552: SAMPLE = 16'ha128;
		3553: SAMPLE = 16'ha14a;
		3554: SAMPLE = 16'ha16c;
		3555: SAMPLE = 16'ha18e;
		3556: SAMPLE = 16'ha1af;
		3557: SAMPLE = 16'ha1d2;
		3558: SAMPLE = 16'ha1f4;
		3559: SAMPLE = 16'ha216;
		3560: SAMPLE = 16'ha238;
		3561: SAMPLE = 16'ha25a;
		3562: SAMPLE = 16'ha27c;
		3563: SAMPLE = 16'ha29f;
		3564: SAMPLE = 16'ha2c1;
		3565: SAMPLE = 16'ha2e4;
		3566: SAMPLE = 16'ha306;
		3567: SAMPLE = 16'ha329;
		3568: SAMPLE = 16'ha34b;
		3569: SAMPLE = 16'ha36e;
		3570: SAMPLE = 16'ha391;
		3571: SAMPLE = 16'ha3b4;
		3572: SAMPLE = 16'ha3d6;
		3573: SAMPLE = 16'ha3f9;
		3574: SAMPLE = 16'ha41c;
		3575: SAMPLE = 16'ha43f;
		3576: SAMPLE = 16'ha462;
		3577: SAMPLE = 16'ha486;
		3578: SAMPLE = 16'ha4a9;
		3579: SAMPLE = 16'ha4cc;
		3580: SAMPLE = 16'ha4ef;
		3581: SAMPLE = 16'ha513;
		3582: SAMPLE = 16'ha536;
		3583: SAMPLE = 16'ha55a;
		3584: SAMPLE = 16'ha57d;
		3585: SAMPLE = 16'ha5a1;
		3586: SAMPLE = 16'ha5c4;
		3587: SAMPLE = 16'ha5e8;
		3588: SAMPLE = 16'ha60c;
		3589: SAMPLE = 16'ha62f;
		3590: SAMPLE = 16'ha653;
		3591: SAMPLE = 16'ha677;
		3592: SAMPLE = 16'ha69b;
		3593: SAMPLE = 16'ha6bf;
		3594: SAMPLE = 16'ha6e3;
		3595: SAMPLE = 16'ha707;
		3596: SAMPLE = 16'ha72b;
		3597: SAMPLE = 16'ha750;
		3598: SAMPLE = 16'ha774;
		3599: SAMPLE = 16'ha798;
		3600: SAMPLE = 16'ha7bd;
		3601: SAMPLE = 16'ha7e1;
		3602: SAMPLE = 16'ha806;
		3603: SAMPLE = 16'ha82a;
		3604: SAMPLE = 16'ha84f;
		3605: SAMPLE = 16'ha873;
		3606: SAMPLE = 16'ha898;
		3607: SAMPLE = 16'ha8bd;
		3608: SAMPLE = 16'ha8e2;
		3609: SAMPLE = 16'ha906;
		3610: SAMPLE = 16'ha92b;
		3611: SAMPLE = 16'ha950;
		3612: SAMPLE = 16'ha975;
		3613: SAMPLE = 16'ha99a;
		3614: SAMPLE = 16'ha9bf;
		3615: SAMPLE = 16'ha9e5;
		3616: SAMPLE = 16'haa0a;
		3617: SAMPLE = 16'haa2f;
		3618: SAMPLE = 16'haa54;
		3619: SAMPLE = 16'haa7a;
		3620: SAMPLE = 16'haa9f;
		3621: SAMPLE = 16'haac5;
		3622: SAMPLE = 16'haaea;
		3623: SAMPLE = 16'hab10;
		3624: SAMPLE = 16'hab35;
		3625: SAMPLE = 16'hab5b;
		3626: SAMPLE = 16'hab81;
		3627: SAMPLE = 16'haba7;
		3628: SAMPLE = 16'habcc;
		3629: SAMPLE = 16'habf2;
		3630: SAMPLE = 16'hac18;
		3631: SAMPLE = 16'hac3e;
		3632: SAMPLE = 16'hac64;
		3633: SAMPLE = 16'hac8a;
		3634: SAMPLE = 16'hacb1;
		3635: SAMPLE = 16'hacd7;
		3636: SAMPLE = 16'hacfd;
		3637: SAMPLE = 16'had23;
		3638: SAMPLE = 16'had4a;
		3639: SAMPLE = 16'had70;
		3640: SAMPLE = 16'had96;
		3641: SAMPLE = 16'hadbd;
		3642: SAMPLE = 16'hade3;
		3643: SAMPLE = 16'hae0a;
		3644: SAMPLE = 16'hae31;
		3645: SAMPLE = 16'hae57;
		3646: SAMPLE = 16'hae7e;
		3647: SAMPLE = 16'haea5;
		3648: SAMPLE = 16'haecc;
		3649: SAMPLE = 16'haef3;
		3650: SAMPLE = 16'haf1a;
		3651: SAMPLE = 16'haf40;
		3652: SAMPLE = 16'haf68;
		3653: SAMPLE = 16'haf8f;
		3654: SAMPLE = 16'hafb6;
		3655: SAMPLE = 16'hafdd;
		3656: SAMPLE = 16'hb004;
		3657: SAMPLE = 16'hb02b;
		3658: SAMPLE = 16'hb053;
		3659: SAMPLE = 16'hb07a;
		3660: SAMPLE = 16'hb0a1;
		3661: SAMPLE = 16'hb0c9;
		3662: SAMPLE = 16'hb0f0;
		3663: SAMPLE = 16'hb118;
		3664: SAMPLE = 16'hb140;
		3665: SAMPLE = 16'hb167;
		3666: SAMPLE = 16'hb18f;
		3667: SAMPLE = 16'hb1b7;
		3668: SAMPLE = 16'hb1de;
		3669: SAMPLE = 16'hb206;
		3670: SAMPLE = 16'hb22e;
		3671: SAMPLE = 16'hb256;
		3672: SAMPLE = 16'hb27e;
		3673: SAMPLE = 16'hb2a6;
		3674: SAMPLE = 16'hb2ce;
		3675: SAMPLE = 16'hb2f6;
		3676: SAMPLE = 16'hb31e;
		3677: SAMPLE = 16'hb347;
		3678: SAMPLE = 16'hb36f;
		3679: SAMPLE = 16'hb397;
		3680: SAMPLE = 16'hb3c0;
		3681: SAMPLE = 16'hb3e8;
		3682: SAMPLE = 16'hb410;
		3683: SAMPLE = 16'hb439;
		3684: SAMPLE = 16'hb461;
		3685: SAMPLE = 16'hb48a;
		3686: SAMPLE = 16'hb4b3;
		3687: SAMPLE = 16'hb4db;
		3688: SAMPLE = 16'hb504;
		3689: SAMPLE = 16'hb52d;
		3690: SAMPLE = 16'hb556;
		3691: SAMPLE = 16'hb57e;
		3692: SAMPLE = 16'hb5a7;
		3693: SAMPLE = 16'hb5d0;
		3694: SAMPLE = 16'hb5f9;
		3695: SAMPLE = 16'hb622;
		3696: SAMPLE = 16'hb64b;
		3697: SAMPLE = 16'hb675;
		3698: SAMPLE = 16'hb69e;
		3699: SAMPLE = 16'hb6c7;
		3700: SAMPLE = 16'hb6f0;
		3701: SAMPLE = 16'hb719;
		3702: SAMPLE = 16'hb743;
		3703: SAMPLE = 16'hb76c;
		3704: SAMPLE = 16'hb796;
		3705: SAMPLE = 16'hb7bf;
		3706: SAMPLE = 16'hb7e9;
		3707: SAMPLE = 16'hb812;
		3708: SAMPLE = 16'hb83c;
		3709: SAMPLE = 16'hb865;
		3710: SAMPLE = 16'hb88f;
		3711: SAMPLE = 16'hb8b9;
		3712: SAMPLE = 16'hb8e3;
		3713: SAMPLE = 16'hb90c;
		3714: SAMPLE = 16'hb936;
		3715: SAMPLE = 16'hb960;
		3716: SAMPLE = 16'hb98a;
		3717: SAMPLE = 16'hb9b4;
		3718: SAMPLE = 16'hb9de;
		3719: SAMPLE = 16'hba08;
		3720: SAMPLE = 16'hba32;
		3721: SAMPLE = 16'hba5c;
		3722: SAMPLE = 16'hba87;
		3723: SAMPLE = 16'hbab1;
		3724: SAMPLE = 16'hbadb;
		3725: SAMPLE = 16'hbb05;
		3726: SAMPLE = 16'hbb30;
		3727: SAMPLE = 16'hbb5a;
		3728: SAMPLE = 16'hbb85;
		3729: SAMPLE = 16'hbbaf;
		3730: SAMPLE = 16'hbbda;
		3731: SAMPLE = 16'hbc04;
		3732: SAMPLE = 16'hbc2f;
		3733: SAMPLE = 16'hbc5a;
		3734: SAMPLE = 16'hbc84;
		3735: SAMPLE = 16'hbcaf;
		3736: SAMPLE = 16'hbcda;
		3737: SAMPLE = 16'hbd05;
		3738: SAMPLE = 16'hbd2f;
		3739: SAMPLE = 16'hbd5a;
		3740: SAMPLE = 16'hbd85;
		3741: SAMPLE = 16'hbdb0;
		3742: SAMPLE = 16'hbddb;
		3743: SAMPLE = 16'hbe06;
		3744: SAMPLE = 16'hbe31;
		3745: SAMPLE = 16'hbe5d;
		3746: SAMPLE = 16'hbe88;
		3747: SAMPLE = 16'hbeb3;
		3748: SAMPLE = 16'hbede;
		3749: SAMPLE = 16'hbf09;
		3750: SAMPLE = 16'hbf35;
		3751: SAMPLE = 16'hbf60;
		3752: SAMPLE = 16'hbf8c;
		3753: SAMPLE = 16'hbfb7;
		3754: SAMPLE = 16'hbfe2;
		3755: SAMPLE = 16'hc00e;
		3756: SAMPLE = 16'hc03a;
		3757: SAMPLE = 16'hc065;
		3758: SAMPLE = 16'hc091;
		3759: SAMPLE = 16'hc0bc;
		3760: SAMPLE = 16'hc0e8;
		3761: SAMPLE = 16'hc114;
		3762: SAMPLE = 16'hc140;
		3763: SAMPLE = 16'hc16c;
		3764: SAMPLE = 16'hc197;
		3765: SAMPLE = 16'hc1c3;
		3766: SAMPLE = 16'hc1ef;
		3767: SAMPLE = 16'hc21b;
		3768: SAMPLE = 16'hc247;
		3769: SAMPLE = 16'hc273;
		3770: SAMPLE = 16'hc29f;
		3771: SAMPLE = 16'hc2cc;
		3772: SAMPLE = 16'hc2f8;
		3773: SAMPLE = 16'hc324;
		3774: SAMPLE = 16'hc350;
		3775: SAMPLE = 16'hc37c;
		3776: SAMPLE = 16'hc3a9;
		3777: SAMPLE = 16'hc3d5;
		3778: SAMPLE = 16'hc402;
		3779: SAMPLE = 16'hc42e;
		3780: SAMPLE = 16'hc45a;
		3781: SAMPLE = 16'hc487;
		3782: SAMPLE = 16'hc4b3;
		3783: SAMPLE = 16'hc4e0;
		3784: SAMPLE = 16'hc50d;
		3785: SAMPLE = 16'hc539;
		3786: SAMPLE = 16'hc566;
		3787: SAMPLE = 16'hc593;
		3788: SAMPLE = 16'hc5bf;
		3789: SAMPLE = 16'hc5ec;
		3790: SAMPLE = 16'hc619;
		3791: SAMPLE = 16'hc646;
		3792: SAMPLE = 16'hc673;
		3793: SAMPLE = 16'hc6a0;
		3794: SAMPLE = 16'hc6cd;
		3795: SAMPLE = 16'hc6f9;
		3796: SAMPLE = 16'hc727;
		3797: SAMPLE = 16'hc754;
		3798: SAMPLE = 16'hc781;
		3799: SAMPLE = 16'hc7ae;
		3800: SAMPLE = 16'hc7db;
		3801: SAMPLE = 16'hc808;
		3802: SAMPLE = 16'hc835;
		3803: SAMPLE = 16'hc863;
		3804: SAMPLE = 16'hc890;
		3805: SAMPLE = 16'hc8bd;
		3806: SAMPLE = 16'hc8eb;
		3807: SAMPLE = 16'hc918;
		3808: SAMPLE = 16'hc945;
		3809: SAMPLE = 16'hc973;
		3810: SAMPLE = 16'hc9a0;
		3811: SAMPLE = 16'hc9ce;
		3812: SAMPLE = 16'hc9fb;
		3813: SAMPLE = 16'hca29;
		3814: SAMPLE = 16'hca57;
		3815: SAMPLE = 16'hca84;
		3816: SAMPLE = 16'hcab2;
		3817: SAMPLE = 16'hcae0;
		3818: SAMPLE = 16'hcb0d;
		3819: SAMPLE = 16'hcb3b;
		3820: SAMPLE = 16'hcb69;
		3821: SAMPLE = 16'hcb97;
		3822: SAMPLE = 16'hcbc5;
		3823: SAMPLE = 16'hcbf3;
		3824: SAMPLE = 16'hcc21;
		3825: SAMPLE = 16'hcc4f;
		3826: SAMPLE = 16'hcc7d;
		3827: SAMPLE = 16'hccab;
		3828: SAMPLE = 16'hccd9;
		3829: SAMPLE = 16'hcd07;
		3830: SAMPLE = 16'hcd35;
		3831: SAMPLE = 16'hcd63;
		3832: SAMPLE = 16'hcd91;
		3833: SAMPLE = 16'hcdbf;
		3834: SAMPLE = 16'hcdee;
		3835: SAMPLE = 16'hce1c;
		3836: SAMPLE = 16'hce4a;
		3837: SAMPLE = 16'hce79;
		3838: SAMPLE = 16'hcea7;
		3839: SAMPLE = 16'hced5;
		3840: SAMPLE = 16'hcf04;
		3841: SAMPLE = 16'hcf32;
		3842: SAMPLE = 16'hcf61;
		3843: SAMPLE = 16'hcf8f;
		3844: SAMPLE = 16'hcfbe;
		3845: SAMPLE = 16'hcfec;
		3846: SAMPLE = 16'hd01b;
		3847: SAMPLE = 16'hd04a;
		3848: SAMPLE = 16'hd078;
		3849: SAMPLE = 16'hd0a7;
		3850: SAMPLE = 16'hd0d6;
		3851: SAMPLE = 16'hd104;
		3852: SAMPLE = 16'hd133;
		3853: SAMPLE = 16'hd162;
		3854: SAMPLE = 16'hd191;
		3855: SAMPLE = 16'hd1c0;
		3856: SAMPLE = 16'hd1ee;
		3857: SAMPLE = 16'hd21d;
		3858: SAMPLE = 16'hd24c;
		3859: SAMPLE = 16'hd27b;
		3860: SAMPLE = 16'hd2aa;
		3861: SAMPLE = 16'hd2d9;
		3862: SAMPLE = 16'hd308;
		3863: SAMPLE = 16'hd337;
		3864: SAMPLE = 16'hd367;
		3865: SAMPLE = 16'hd396;
		3866: SAMPLE = 16'hd3c5;
		3867: SAMPLE = 16'hd3f4;
		3868: SAMPLE = 16'hd423;
		3869: SAMPLE = 16'hd452;
		3870: SAMPLE = 16'hd482;
		3871: SAMPLE = 16'hd4b1;
		3872: SAMPLE = 16'hd4e0;
		3873: SAMPLE = 16'hd510;
		3874: SAMPLE = 16'hd53f;
		3875: SAMPLE = 16'hd56e;
		3876: SAMPLE = 16'hd59e;
		3877: SAMPLE = 16'hd5cd;
		3878: SAMPLE = 16'hd5fd;
		3879: SAMPLE = 16'hd62c;
		3880: SAMPLE = 16'hd65c;
		3881: SAMPLE = 16'hd68b;
		3882: SAMPLE = 16'hd6bb;
		3883: SAMPLE = 16'hd6ea;
		3884: SAMPLE = 16'hd71a;
		3885: SAMPLE = 16'hd74a;
		3886: SAMPLE = 16'hd779;
		3887: SAMPLE = 16'hd7a9;
		3888: SAMPLE = 16'hd7d9;
		3889: SAMPLE = 16'hd809;
		3890: SAMPLE = 16'hd838;
		3891: SAMPLE = 16'hd868;
		3892: SAMPLE = 16'hd898;
		3893: SAMPLE = 16'hd8c8;
		3894: SAMPLE = 16'hd8f8;
		3895: SAMPLE = 16'hd927;
		3896: SAMPLE = 16'hd957;
		3897: SAMPLE = 16'hd987;
		3898: SAMPLE = 16'hd9b7;
		3899: SAMPLE = 16'hd9e7;
		3900: SAMPLE = 16'hda17;
		3901: SAMPLE = 16'hda47;
		3902: SAMPLE = 16'hda77;
		3903: SAMPLE = 16'hdaa7;
		3904: SAMPLE = 16'hdad7;
		3905: SAMPLE = 16'hdb08;
		3906: SAMPLE = 16'hdb38;
		3907: SAMPLE = 16'hdb68;
		3908: SAMPLE = 16'hdb98;
		3909: SAMPLE = 16'hdbc8;
		3910: SAMPLE = 16'hdbf8;
		3911: SAMPLE = 16'hdc29;
		3912: SAMPLE = 16'hdc59;
		3913: SAMPLE = 16'hdc89;
		3914: SAMPLE = 16'hdcba;
		3915: SAMPLE = 16'hdcea;
		3916: SAMPLE = 16'hdd1a;
		3917: SAMPLE = 16'hdd4b;
		3918: SAMPLE = 16'hdd7b;
		3919: SAMPLE = 16'hddab;
		3920: SAMPLE = 16'hdddc;
		3921: SAMPLE = 16'hde0c;
		3922: SAMPLE = 16'hde3d;
		3923: SAMPLE = 16'hde6d;
		3924: SAMPLE = 16'hde9e;
		3925: SAMPLE = 16'hdece;
		3926: SAMPLE = 16'hdeff;
		3927: SAMPLE = 16'hdf2f;
		3928: SAMPLE = 16'hdf60;
		3929: SAMPLE = 16'hdf91;
		3930: SAMPLE = 16'hdfc1;
		3931: SAMPLE = 16'hdff2;
		3932: SAMPLE = 16'he023;
		3933: SAMPLE = 16'he053;
		3934: SAMPLE = 16'he084;
		3935: SAMPLE = 16'he0b5;
		3936: SAMPLE = 16'he0e6;
		3937: SAMPLE = 16'he116;
		3938: SAMPLE = 16'he147;
		3939: SAMPLE = 16'he178;
		3940: SAMPLE = 16'he1a9;
		3941: SAMPLE = 16'he1da;
		3942: SAMPLE = 16'he20a;
		3943: SAMPLE = 16'he23b;
		3944: SAMPLE = 16'he26c;
		3945: SAMPLE = 16'he29d;
		3946: SAMPLE = 16'he2ce;
		3947: SAMPLE = 16'he2ff;
		3948: SAMPLE = 16'he330;
		3949: SAMPLE = 16'he361;
		3950: SAMPLE = 16'he392;
		3951: SAMPLE = 16'he3c3;
		3952: SAMPLE = 16'he3f4;
		3953: SAMPLE = 16'he425;
		3954: SAMPLE = 16'he456;
		3955: SAMPLE = 16'he487;
		3956: SAMPLE = 16'he4b8;
		3957: SAMPLE = 16'he4e9;
		3958: SAMPLE = 16'he51b;
		3959: SAMPLE = 16'he54c;
		3960: SAMPLE = 16'he57d;
		3961: SAMPLE = 16'he5ae;
		3962: SAMPLE = 16'he5df;
		3963: SAMPLE = 16'he610;
		3964: SAMPLE = 16'he642;
		3965: SAMPLE = 16'he673;
		3966: SAMPLE = 16'he6a4;
		3967: SAMPLE = 16'he6d5;
		3968: SAMPLE = 16'he707;
		3969: SAMPLE = 16'he738;
		3970: SAMPLE = 16'he769;
		3971: SAMPLE = 16'he79b;
		3972: SAMPLE = 16'he7cc;
		3973: SAMPLE = 16'he7fd;
		3974: SAMPLE = 16'he82f;
		3975: SAMPLE = 16'he860;
		3976: SAMPLE = 16'he892;
		3977: SAMPLE = 16'he8c3;
		3978: SAMPLE = 16'he8f5;
		3979: SAMPLE = 16'he926;
		3980: SAMPLE = 16'he957;
		3981: SAMPLE = 16'he989;
		3982: SAMPLE = 16'he9ba;
		3983: SAMPLE = 16'he9ec;
		3984: SAMPLE = 16'hea1d;
		3985: SAMPLE = 16'hea4f;
		3986: SAMPLE = 16'hea80;
		3987: SAMPLE = 16'heab2;
		3988: SAMPLE = 16'heae4;
		3989: SAMPLE = 16'heb15;
		3990: SAMPLE = 16'heb47;
		3991: SAMPLE = 16'heb78;
		3992: SAMPLE = 16'hebaa;
		3993: SAMPLE = 16'hebdc;
		3994: SAMPLE = 16'hec0d;
		3995: SAMPLE = 16'hec3f;
		3996: SAMPLE = 16'hec71;
		3997: SAMPLE = 16'heca2;
		3998: SAMPLE = 16'hecd4;
		3999: SAMPLE = 16'hed06;
		4000: SAMPLE = 16'hed37;
		4001: SAMPLE = 16'hed69;
		4002: SAMPLE = 16'hed9b;
		4003: SAMPLE = 16'hedcd;
		4004: SAMPLE = 16'hedfe;
		4005: SAMPLE = 16'hee30;
		4006: SAMPLE = 16'hee62;
		4007: SAMPLE = 16'hee94;
		4008: SAMPLE = 16'heec6;
		4009: SAMPLE = 16'heef7;
		4010: SAMPLE = 16'hef29;
		4011: SAMPLE = 16'hef5b;
		4012: SAMPLE = 16'hef8d;
		4013: SAMPLE = 16'hefbf;
		4014: SAMPLE = 16'heff1;
		4015: SAMPLE = 16'hf022;
		4016: SAMPLE = 16'hf054;
		4017: SAMPLE = 16'hf086;
		4018: SAMPLE = 16'hf0b8;
		4019: SAMPLE = 16'hf0ea;
		4020: SAMPLE = 16'hf11c;
		4021: SAMPLE = 16'hf14e;
		4022: SAMPLE = 16'hf180;
		4023: SAMPLE = 16'hf1b2;
		4024: SAMPLE = 16'hf1e4;
		4025: SAMPLE = 16'hf216;
		4026: SAMPLE = 16'hf248;
		4027: SAMPLE = 16'hf27a;
		4028: SAMPLE = 16'hf2ac;
		4029: SAMPLE = 16'hf2de;
		4030: SAMPLE = 16'hf310;
		4031: SAMPLE = 16'hf342;
		4032: SAMPLE = 16'hf374;
		4033: SAMPLE = 16'hf3a6;
		4034: SAMPLE = 16'hf3d8;
		4035: SAMPLE = 16'hf40a;
		4036: SAMPLE = 16'hf43c;
		4037: SAMPLE = 16'hf46e;
		4038: SAMPLE = 16'hf4a0;
		4039: SAMPLE = 16'hf4d2;
		4040: SAMPLE = 16'hf504;
		4041: SAMPLE = 16'hf536;
		4042: SAMPLE = 16'hf568;
		4043: SAMPLE = 16'hf59a;
		4044: SAMPLE = 16'hf5cc;
		4045: SAMPLE = 16'hf5ff;
		4046: SAMPLE = 16'hf631;
		4047: SAMPLE = 16'hf663;
		4048: SAMPLE = 16'hf695;
		4049: SAMPLE = 16'hf6c7;
		4050: SAMPLE = 16'hf6f9;
		4051: SAMPLE = 16'hf72b;
		4052: SAMPLE = 16'hf75d;
		4053: SAMPLE = 16'hf790;
		4054: SAMPLE = 16'hf7c2;
		4055: SAMPLE = 16'hf7f4;
		4056: SAMPLE = 16'hf826;
		4057: SAMPLE = 16'hf858;
		4058: SAMPLE = 16'hf88a;
		4059: SAMPLE = 16'hf8bd;
		4060: SAMPLE = 16'hf8ef;
		4061: SAMPLE = 16'hf921;
		4062: SAMPLE = 16'hf953;
		4063: SAMPLE = 16'hf985;
		4064: SAMPLE = 16'hf9b8;
		4065: SAMPLE = 16'hf9ea;
		4066: SAMPLE = 16'hfa1c;
		4067: SAMPLE = 16'hfa4e;
		4068: SAMPLE = 16'hfa80;
		4069: SAMPLE = 16'hfab3;
		4070: SAMPLE = 16'hfae5;
		4071: SAMPLE = 16'hfb17;
		4072: SAMPLE = 16'hfb49;
		4073: SAMPLE = 16'hfb7c;
		4074: SAMPLE = 16'hfbae;
		4075: SAMPLE = 16'hfbe0;
		4076: SAMPLE = 16'hfc12;
		4077: SAMPLE = 16'hfc45;
		4078: SAMPLE = 16'hfc77;
		4079: SAMPLE = 16'hfca9;
		4080: SAMPLE = 16'hfcdb;
		4081: SAMPLE = 16'hfd0e;
		4082: SAMPLE = 16'hfd40;
		4083: SAMPLE = 16'hfd72;
		4084: SAMPLE = 16'hfda4;
		4085: SAMPLE = 16'hfdd7;
		4086: SAMPLE = 16'hfe09;
		4087: SAMPLE = 16'hfe3b;
		4088: SAMPLE = 16'hfe6d;
		4089: SAMPLE = 16'hfea0;
		4090: SAMPLE = 16'hfed2;
		4091: SAMPLE = 16'hff04;
		4092: SAMPLE = 16'hff36;
		4093: SAMPLE = 16'hff69;
		4094: SAMPLE = 16'hff9b;
		4095: SAMPLE = 16'hffcd;
	endcase

end

endmodule
