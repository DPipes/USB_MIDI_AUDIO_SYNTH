module f_table(input logic [6:0] KEY,
					output logic [23:0] F
					);

always_comb begin
	case (KEY) 
		12: F = 24'h184c;
		13: F = 24'h19be;
		14: F = 24'h1b46;
		15: F = 24'h1ce5;
		16: F = 24'h1e9d;
		17: F = 24'h206f;
		18: F = 24'h225d;
		19: F = 24'h2468;
		20: F = 24'h2692;
		21: F = 24'h28dd;
		22: F = 24'h2b4b;
		23: F = 24'h2dde;
		24: F = 24'h3099;
		25: F = 24'h337c;
		26: F = 24'h368c;
		27: F = 24'h39cb;
		28: F = 24'h3d3a;
		29: F = 24'h40de;
		30: F = 24'h44ba;
		31: F = 24'h48d0;
		32: F = 24'h4d24;
		33: F = 24'h51bb;
		34: F = 24'h5697;
		35: F = 24'h5bbd;
		36: F = 24'h6131;
		37: F = 24'h66f9;
		38: F = 24'h6d18;
		39: F = 24'h7395;
		40: F = 24'h7a75;
		41: F = 24'h81bd;
		42: F = 24'h8974;
		43: F = 24'h91a0;
		44: F = 24'h9a49;
		45: F = 24'ha375;
		46: F = 24'had2d;
		47: F = 24'hb77a;
		48: F = 24'hc263;
		49: F = 24'hcdf2;
		50: F = 24'hda31;
		51: F = 24'he72a;
		52: F = 24'hf4e9;
		53: F = 24'h10379;
		54: F = 24'h112e7;
		55: F = 24'h12340;
		56: F = 24'h13491;
		57: F = 24'h146eb;
		58: F = 24'h15a5b;
		59: F = 24'h16ef3;
		60: F = 24'h184c5;
		61: F = 24'h19be3;
		62: F = 24'h1b461;
		63: F = 24'h1ce54;
		64: F = 24'h1e9d2;
		65: F = 24'h206f2;
		66: F = 24'h225ce;
		67: F = 24'h24680;
		68: F = 24'h26923;
		69: F = 24'h28dd5;
		70: F = 24'h2b4b6;
		71: F = 24'h2dde7;
		72: F = 24'h3098b;
		73: F = 24'h337c7;
		74: F = 24'h368c3;
		75: F = 24'h39ca8;
		76: F = 24'h3d3a4;
		77: F = 24'h40de5;
		78: F = 24'h44b9c;
		79: F = 24'h48cff;
		80: F = 24'h4d245;
		81: F = 24'h51baa;
		82: F = 24'h5696c;
		83: F = 24'h5bbce;
		84: F = 24'h61315;
		85: F = 24'h66f8e;
		86: F = 24'h6d186;
		87: F = 24'h73951;
		88: F = 24'h7a748;
		89: F = 24'h81bca;
		90: F = 24'h89738;
		91: F = 24'h919fe;
		92: F = 24'h9a48b;
		93: F = 24'ha3754;
		94: F = 24'had2d8;
		95: F = 24'hb779b;
		96: F = 24'hc262b;
		97: F = 24'hcdf1b;
		98: F = 24'hda30b;
		99: F = 24'he72a2;
		100: F = 24'hf4e90;
		101: F = 24'h103793;
		102: F = 24'h112e71;
		103: F = 24'h1233fc;
		104: F = 24'h134915;
		105: F = 24'h146ea8;
		106: F = 24'h15a5b0;
		107: F = 24'h16ef36;
		108: F = 24'h184c55;
		109: F = 24'h19be37;
		110: F = 24'h1b4617;
		111: F = 24'h1ce544;
		112: F = 24'h1e9d21;
		113: F = 24'h206f26;
		114: F = 24'h225ce1;
		115: F = 24'h2467f8;
		116: F = 24'h26922a;
		117: F = 24'h28dd50;
		118: F = 24'h2b4b60;
		119: F = 24'h2dde6d;
		default: F = 24'h0;
	endcase
end

endmodule
